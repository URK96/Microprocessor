XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����p�E�ß�R'[���]��d��u{�~G�܂���',�J.�b�xY�F��Pg�^#x������p����}p�!�hm	~D1���P�R���<%��>�ľ��ѥ�F��E"\�	}Z�m	��w��D:���x��b�]�$+�<�xV�	H x����b��ZR*B:{N�������M���ӮvKVJ)�<��1��OU�N��f��X�Ȝ�"F,�.��&�'3%��p�x$�Bά��{��%��y#%�	О�$��\�X�V87��5���=��=�sƹ-�G�	Q2ߩօ��R�D��UKW�* �{�����)@D����&V<5�X�.���վ�샧������Bb*Nv;(��,����i8G��o��m_-�]���R�v�� �v��\�"!{?�w����y�+��Uu��flz��]+�&���8�ɲc.�$�M?���K�,��q�g�LƘ_�:�&J��q�'����Ͼ���n�-.Ҹ&�$[���VS�n� iw�W`��'*�7���'�bO,�ۇ~��k��$�Ǆꭀhj߲a$I9�ޖy��#wgz��F���������$y�:�Dhz� 2�Q8�"��}��s@U���%�;�W�V��RTey����=w� ��hA�~
�f�<Q��	N>��d�k����ΦΡ�d�9�����zD���6��sQ*l�
�6}�^7Gdn��Y��B�/�T����-K��%q����[�taJ(Ĳa �XlxVHYEB    152b     580,��z�X�Ku�B�r���h;@!8N��OS��AU���ߕz��M��� Ҽy���l�v�V��"���2O`����~:$(����b'�AV:���Ǌ�"0z$D܇D�4!S�,�'��j.�̘|��G�]eg�z�}��Z�W�?�$�fd�8�i�w`k !L��j�留��G���z���^Ք�hͱn���
AAW/�p[��B8���XpѶ�a"�r��*�>�#���P�.T5�ӉA%�B�6��8�=0�K��:A�eȎq��>�]X���=-���zb"����	��4.Yot��أT����)MQ�x��A�7pP��:s���Z�_�R��.���BA���l��l��G���J��*��eY =�r�P{�ZqˢŒI��
EJ��v��~��E��Ȇ�50NZz���-���G?����3�h:{�Hӄ��O�?��wX@Tw��ݞ4�ƹc}��æ<h��J����5K��?��^�K\;��Zx_!�J�����J(,���#�"6��Q��lT
0Ӹ��~*|�{HF�M�F�p�Oməo�O2�	ƛA/c���%�+j�)� ��8z~��l7BX�4�~��3�v����2��Қ�\�\}B����q �y1c��r��m���r
`��DYK�7��i�(��,�5ȶ�C6����a��ù$�E�PˋN��"��]_�э����[��S��$�*oI�e��^^�����Ϟ�şv�8i�j�AB=>@�rk���"	�����ط����Ѫ��?�E���FUҨKf}0��)�=��~��Mv��i z@#<��<a�b�w R2uS�����jp��>Yؐ�!�t�^��?�0��q[
=�� ��.F��
w0�Rw^Z�J^���aa���s��%���:��`~J:
����� �S�N�>&�N;c�Ap�	��������|S�w$�h��d�	+N�Ƒ���J����A�A�3ĩ2 9k��n�Xx�"�FD� Q���1�	���1��,�Ыk�n��X?��a�ytj��#A��N�ADW��H�2�UT��k��B�m R�=Z�%-Bf�d�)R�:���ed	6Nn_��}с�^�-_�l�Y�yV.]vk���}8���Gm�� ��������>n��E ,���"����ug4�b�8TQ�J�y�$��t�m�˭���u�����d�E����T{��bD߂/f:��\�n���ߤ�Xc�{y��F���NR�Y�C��= ���
�΁QYL^��W��1������9����'}�C��P�]���Χ��QK��L�'�>��j���WkH�pܰ���Q�,�5	�}ӱ��?������T	���5���oo