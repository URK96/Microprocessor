XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����Sh*�Q�!�.d_v�pT|�T]gr\t�[{�Q�x9�{�9�V�_*�R@)S���τ�=f��Ka�X,�t���9T����A3�Q~���me��c�M��*�"F�-bU(K��~������yJ�+���+-���0E�4��������U����Z����0�P�y�r���x_4��0��Fw��"��Eu�«\q�.4�I0��ή�m.�}[\~:{�3��D�Rs��H�4V˸�s�v[�c6�F���|��jF�6t�(ɏ�f�~]hs(�ץ�}��;�w}5أ��F��,���m�7�-%Z�*Y��bSS�K�K�����[GQk���"��-H��T!�­�W�U�$9P����ÀF|��x���~�^�h��L�*/��o�`(�ћD� �keԡ6l��*��#���w-u�����,�fvP���;�J�W��\xJ������`#�)��Wi9ͦ+�h�f��
Y����	����I(���p���E�!�5�նK�U����o��LF7���F6Ԫh���x�N]�j~ȵ���F+Ԡ����E݈�R��9k}�8֖�d+Fa8k%��� �V@v�.;fC^���a����H$#�b	w�d r�WP�Ǫs��T�>��0ճZy"}��)	�3ktPl����Vk�v��f=�>���ͦx,����ׂ������"x�P�d���-,69�-���q6��6L����/k�2K��ns�1���rBXlxVHYEB    cc3b    16b03�w�����/3�D���2�����O����������\.�}	z���=����eAl�T��'V]��?�ym�Z(���&8�%ä|i���s��>]Q;@@�H"���iq��f�H��=�*��k��ݪ��]������ L!�����IO�l�6�[�TE�ĲUGm)F�0-�B�ɏH�|K���.Q�u�c��K:U��i�L��<|�]�Ռ�&�%m��$Q�6j��Ȕ��I@���p(�?�
�FȀ������%4����ҿ��Z/�.���Z������N~+Sĥ[��⭜!�'�����E)%މ;��l�T��}��0t�Ds�m򫟮�OЊL���vf-��5pz�)��^4
yK-r�>�6��<݀��<��	�*��} ��$�}���5�Xl�����jDI�Þ������ST
zT�v໖%?	���q-�dJp'S�z�K�K?<n$��2}fF�ҷ�	���cO�,D�8�UX�'I�w���Dm�6&�L��1o!��	RVS�#!��&C|�YeL2�W3�5�k[Ή�с`(��"��	~�Tҫz�K"L�^����J������1�M����D���4ڔ�	Ie�@�����Cg�1��4Ϧ9yC����B�og�&����|���`H�Swċ���
V&��ٸ�kri\��mx���TW��nrs�߾0G!�áQ���{ƈ��ϔ�a��w�Q�����U�7�I�F>�����+uGI�z_���4}�d����ЮX��%xiYx�hE�ڋ��.�sIX�H�.T���?�;U�J�S=�����р�i2#��nc��g��tu��Z
h���wė%d�9z��&J���c/��Ce��]t��j��Wq���X7$[�#@���oUW����`u�Z�v\h�P��xm�I���"��s�R�+��D��j�>({��/�`����(8ĸ���E����p�Z�g��8e�Rؐ��~P�\ۋ=��Z(��g�a� ��O@�WC�� f;L�c���.��'��Vʙ�K'
Ϋ�Dx���<��OjK����<k��HG�N��Q��e^k$�ʬ&V.��i�b!UӀ5������@����)O�����+�LwU�}�4]Q������?��;����߽�A�,��F���٢�Nⷫ�z�-?k=���9D��0��{�v�
%*?�.8z����'��
Y�q���_R�V�8 ZiO��rx�z���~u�\��Md�m�_���ἡ�9�>����{� ��&mz��K�J;vU&]Bܵ�%�mq�Sf�8�Jڊ�L�̈�Q��m�Nr�� p�r>Jˑ�-zQ�]�W����F�ukmݞ1�Ƒeh/κv)9J_��7�.�����׌Ҵ���FC��?P���x����?�
a��Zy��Wi0��)������C�}���$�^u@��`��8�K1/�m���Q��a*)j��`"˩���?��k�u4�\�v�c��(�&�LV�~-<b*�u1����V����Hw��&���������.p�����6b� �;��΀;�R8|7��"��{����5���On��W�wm����R$W4���UK��_�x�΅_���{e�0/�R3^K��p�"����;�֎��;�X!���`u��_�37�*�j6d�A��I��~@�5��0cKuj{��)��})Hz��g$ȸ�0u����)ܬ��,��&{+�V���
�ɛ��OLD���E`��?)�n(:����fv/��ϊ��Q9Z ��J&���"���met��ε�7���H���*%	�~K�/��hCEiXw�O9H��~[�l�����>��n|��4�1��c�H��g���$�
�g�t�+�QR!x���p��Id��nS��R��'�V�v���U������$��^�5V����Y�]����b�q�C�����7��BE~T��`���j�_ !;$s�Mm�ў`�Ӻٺ��ߐ�k�	��s0�r�z��Y%�҇�]>A^:�e ??�k�� Ԙ>
�`*��<��X2�'��(�q�٩\�'ɍ^�����%�i�g@Ii�QJbM|$�E�ҿZ�dC7w�}*��%|�t*Q�W�Ybi���2<n��7{Ai��iQ�0�d�A��zW�j�������@ϣ<qv��0%�N^�����e����ɷw[O[�3�.j�ݿX�ĜX�Q[�6ba2%��җ���V]R D��eL������eʞ bޭ�0.ݎ�ܰ���=mO���n�y��O(;x���J�>\�\4l�ݩ�KT��@�&PVNC��#�\�g��(w%ގ�}���#��Ik�+
s�)�+bw[GG�)�*��a�IYB��<!QP�L���,"�t��^�ٵ��+�ɋ�A�Ig
�Y �u���!G��G�A�X ��i�+���i&�6���`��&�/�Ow�uڞ�����H�!^MV5�E���~�.%;��+.}��n_4�{v�$��L�pƶZyJ���s �mO'(�|� V�~�Ub�[,��*�"�z�ƹQ��E��2YdY�cS�*����rDh�1F�b�F-��Ԧ��{a�ЫՐ@���S�<%��ψ���=����{�)6�p�=oǷv��u�-������)-�Y��N�I�$h���D��7��ߥ�KvuY�`5��Ӆ�5YA;����?�F{���@�g��m�!ok�"i������	eM���wC����1jyj��7
�;�����b�R&��VFä��'o>c4�>�
�E��VV`�: s`��F�CQz+l�Y)>X�eP��N{�R�7�Z�8��zF�]�(@���:(hL�_wK��!�u`}����(�k�˕��v5��"�|�\V����ح��̩�����1.�Nɺ����Wv��o��p�Z/��o8�$a�DV����Q>8��t�D��)7�f�4�!�mį���(9#��m14��9_��qql��n�1r\��B�q�!9���W�cF�G���(���z~� �pȔP(���F&,S�j�p��űb��$�OV�+d��R�w��*�.*���e׸�)����')v���tɱ�C���?� ���B����m��4�m��;b��#BÅ�'�(�~�ίѓ)t�o�_���D�������#�����S\��h��v�L�]�v�����I�׮��\�0���$�;+G��M����t.vv�\(��Uư�����0�~ᑬU�$�����F�"�S�fA;'��h�C )�Ax��7튎�M:5��ל<`)ӽ����,x�cf�uaT?`'�W"�Ǩ����Hsi{�����.��ar.�����	�^'��!������A�±�,�0{��dL���<Q�=����ߧ�DR�Q��:G����gD�g�k��ɰ�<0Dk�A��e�{s�u��<��ǩ� ���y�ZG=�cy#�O�=,X
����=��"�'35 ��_?TU������M���XdDC�![��}�lS�ĺQb�B:j�L��)u�0�	�i�N���ӊ�Sa留�L��e�Bm�{1Z-���SC�C��k�-6����sQ���2��6�&�>����V���`'�UN\?��g�M7�6E��~2"�wA�I�:�'�iz�#�ڛ�8s�"z����(�PE0���%C�]ۙ����w��գ:DLg����G�er�	�װ���~���~>R+8FEe& ��1�j���I�HD&?�(��3n�{4��FG����4��RQ��P�^ܹ�(*�Y�����9�e����v�:��৮����Խi����bҟ����ڜ���Mu��ފ���렏~���0��X�rӪ'�Y�U�����;������a��=�snW� ���v�������t�z	l�r�_F��e�=�}���rM�"�4r�z	��AT�tk�����ɽ'��
(/�J}�6>����%}FO\H�����Jr	�=syC
���>����������;ZsE������)b���W`�5�;|�I�X���6_h,�D�G��5�]-��me��kJa!���O�-q)~H݄�P���Q5�����<�_� ���q�6hx�{<}3[��}����^�GWii�E��A*9f�6�2O;�����xy�8�]a�>£�B]Ug��EK{e�"�:*� �M�-Ϧ�Z0����wξt"�zt�4x�a������V_�Yb0�e�������O�Pn|I��PW��'sb�j�"%�Tҁ@���N��R܉��2��"!��y 5Lt����?��U���&��jI�`ޡ��
�z�2ȹ.����^P��ԭѼE�=��$�r�68��O�����n9+r7q��l��kO�l�K.$ĝ��`zS��҄�a��`�nt!� &]°�JF�LY���I�Gm0�CH��p���?�域�* kO�w���֫A�̪Qp��y��@pڀ'XNȕz�����^���$��6?>�[�Q�H�)=Cp��� ����Xa�S���t~zB����d}��~^&e&q���� �S�M���E�4����W(F!8��A��$S:�ˤ;|�:�Dm�\;4D#Wx�ki/�<��,Qw��(żQ9|�t۶OY(���N�;��ẍ�~5�E*�¿6I7�2F.�ͩ�*^��<�α��Ӡ]}�_�����������}(WN��
,Go��>��l��WM����sR���ߚ��^ �9Ω��]�p"-���M��ֈ)n�(���(m7��1I��q5e��~�P�~)�L�.m��D-�hR�G4wZ	��:��F�ɉ�CZIs��GS�p*8Q����e����F}�!�J~^�)��g"g��wL*񲡵���C&����nl�ۀ��s.�.!�k
��՞��M7~�j�T�n�EߪZ�C���~	��L��j/tp�_K�IG�ufK�����)�>&��@��7B�q�t���ŋjڳ�R d���)Ѵ���%�ԯh3���,��(%�zS�|�!  D�&D�\B�QGo�'ms*֬'���Y�;��E�m�-TQ��}������_!��"�8�z>|�����l�M�m�����e]�=,��h��u�������$��9�D[�d�����*0Pf�y���C�b�Z�2�~+����ō6@%9}��?�~�-8kF��>oN�46Ǻ��VM�5��-�g��&>����L����s8D���]�tْ_����I���[��YJ�.6�;�CS��k8��>�6�z�\r�l�d2�E���-�}Ah������pZ���r ���w���r�L��	��6u�K掔:a��ar�m��S-�L�.u�^e�ZDQ�[�@�G���k�Ю1Y	���d�Z@6�F�3'eH4j�񍃀��bZ~U��x�Hd��p�E-�8��o/���Rx����䷼��7�����X	Z0x�Z6\~�u�wj_H�斄{����[1B?p�:%�to63{�u
�|O�p��u��tW]̓YrQ֭���à�)�tC�7i�K��u�W�I�T��`�9�Vq�v�	F�T!���ʐ�I��%���7�٩��%�x���"a�Q���E+�"u|0�5��"�Yb�[����+� )�[�5