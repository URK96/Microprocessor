XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m�aN�����q�W��r�A|�����/䌍�D-S[�M�k5Ұ���)Hc�p���oXq�̤����L1�#߂9#����h=��� -^�M�HM]��y7��[L�~��#�	��VC;�U���>�uJ�	��K��sۿ��A�*�_;٭�<a��j�H�nKB$�F�xe �*�3N�@�^��B�.�<x�% ����ɶbi�]E��R�ez���A��Ɋ��qCO8Z,/�b��@Et���zbs�g�F5㒴
�GeJUo'7g�!�g�ǖޯ�V�����S��B�AԞ��˟���	@�匮T1PL����5;R��+P5(��Vi�P�9����c���I��{�))(�%�7F89{�`|p����`8	>GaG�L���tW�y��/��ͺ�$4krhgQK��ps���.;.V�������w��h�UZ�ʅ��/�$���Y�ȭa�S� ? ��ݵjnb����Щ���F1�Gj���&�K ����^���Xf��5`˱�*K�lf.
�B���^�e��!�;�W
>��e��N�`z� �TC�sHS��qs�RNe����J�\ȑ�oq֖�̠ũ��+NP�y.��o��E���K���?���ۨ��#[t�K�l�	�qCz����p��sm�v ��s�Q;�b��ـ�\��>,:�{(ɖt	b�rvO���m�����@H��]���6��JX�!�{�'��8K��<�rrq?�z�:N2������0��u��茤S�YXlxVHYEB    3a1c     d40Z�bE�;���x��!��}�O�v���)c��[� � ��0;yO��|�R����6��̮55��7�b%Oq%��%�RD�R�2���q��T����;�.�C:dr{��j�w���,�?Xê�/�u�
9X�$����w�v44C�s)��g�u����i�0��e�T��{�S��,�ƙ]~�F,�ݸ7�T���������+�&�7f9�M�
眸b��y��t�F;�A�8k���@��v��+���������X��x����[F��E�e��j��\V%{���E���֏�; D�d�O��p\QCU�E����7)|$��S�!�^�Z�Ec�S��H�K��ǯD��| ).C~h˶s4�|�B;�)`�E%&���%��P�t<o83�X�Qx9�Ř�o�-7$ #d�"��;~���c_}�f��6�gf���6wd���4������i����ɽM��Q�y<���&p�0ƒ}����x9����c�Դ��#P��Z���<LO�V�w&��uX �U���h���f{���p�lKWo���I=��B�m�J�%��� ���)t-���(^?�=�273���Ζ��������b��x�_�!���Bd���[�h0�q��r��2H�z��ޭen��nxp>�F*�X�ke9I��H��*ɱ��^$ʽ��6�;����qʝVzܴ�_j�-��W��$�\�W[W1�a,�F%��d�'�m~Jl�B�e�T�ɰZBNw0v V�ja̧Q��]:](d���o؇��2H�^R����jS���H�k��Y51�ӋƘ+�I�`HN#�*�
��d�Ϛ�%�.\��7�6S����&�ЏN�`�����p���ѯ�p��%u�r_*ؗq���.�<0/��Bh�ր�����A9�\�����<3�˝Zୟ�fW/�A�y�g���;�w�@C���j";
��솋B[���'"vK$�R�D���q��"�n�7��:����j<o�@y� s>��A��i<���K3�)��j�s\�$�E�}�&�
'F�#c� ��~~sD>J�\z�+W(��c?G��8��&��S��*W��Y�͟r���Z��:l�P�KK�G;}��Qџ6O&��6�c^�HD湈`w��}��4>QQcld�q�%喲�(�V�R���%�Er��#է�#ỵ����}�����$�31ߪF-M��R6�P��F�=�w*KR�Ami���jC��F���*q�9�69����jw���&���������^��+�j@2�*"�sR���f�P��ɫ� l�!H��a��2�� ��Z���ç�
g<s���t=r1!JTNbP'{|r��j��+S&\�uG$�i�*��*Cl> >�+[�.hh:׆IvFa��Q��_�D(v��&���d~Ƕ�[�0�w6����a4�xY���0�ƣ��tm O}ܳ��XƳ��nlm�'JJx���U;��>�LE'�u�����#������5�HW9T�:���^���D�Ô�ل�QC�>�d���s��)i�{�Q_	�:��N1��;~e�;��r�0S��7���"�&�/�д�1}�[Y��m�2?L���D������~�>c �I;��NJ���C���W���u�:(9�9�t@u�	��^OT�q/�i�^r�ӱ��"���+��QN4
���(pk���$d���V�vQ g]˷a���+L,�#�(ݢkz����3-�8�A^���b��!YWχ�~�j���\�*Iv�1�`)Gs����{C�%��\�b�ޢZ��]��Δ%,��n(q@���$Е.q�+��v���W(/H�����'=NDD��#-�v��a���_?�)�Cu!��ҌM�G�;�>M`�r���e(Oa�Ҭ�`|��A��E�L�wQ���Q�5�d��v��Gb����-�U\?]55�|{Sq�Օ�H[Դ�Vz�����"Vb=�	.8e�1���他.���ֶ�F�rٟp��4�%�����G��FV�o�.���1;�S���Ǒ���8+��=6����v3�&��鱪;�}��$�>�W���F��D�g�������l�]�v[����q��:�+�q�Ǒ���j���29K��
+%�J��+�'$�pUf���N"��=��_�S�3�����" \���?� 1�Q��t%E�ūTY���z�����nu�� �v�׼�_�a�Rq/����i7ǖiׁ��^bچ�6Xv�����૒��0.v��_o(8?�kSA�7#3�Q~�e��Yu�f�x�_m�Jm�.�\��ߒ���؆Y���6:%٧Z��-2�*y+�0ݙ���6��g�=��0�F�W��y�G��t4�܍�"�9a5���͖G��Hx���-�Y�,�L�(��xdY/��G�<W����)���Tr7*k�+v�탰�/�f<8�3O963��HyJ#�����vSU�N� �G~��;�����b��٢��O�BtY�#ң�^Ξ53��j'thΪ�i�d`��hu�1ag6u-3F�	H�U�{]��u����}æ���M��%�ֈպ�OI�0ʁ��Hϋ� ��7n8� >u\H)�TTE_�-� o+ѥ�B�n��.�ӈƃ4d�8�+u!kf�~�˱T/��H�CS���<+U�o7(�M���O���H����{��3�m�G"��j��#D��^����P�S�RA��;�
��]��[��4BX v|D�v=r-�>��M���л����l�{�Zݞ�)���6�9�D��W2�R;9�4fu� F�KN��ˬ��-�N\���?ŉ�S>��6��{z��K������-à��N�O*`�Es��GӇ�hF��}�Ҵ�yxMv��D��R>�b=`��$.�L4�x�C��$�%�KE)�f=6+{����_!���F_��@(�%"���z>��=�,�Q,)x�Ϗ��+;��!FN��ۄ}�;e�$ԜW��m:�j�q����y|����?lX�R[m��i"x]E����M���yR�2]4C�<J�߭8�]!�YrO.9���#�M�=�	���
̖u5�f����[0i�:۩���ʈ�M�H��2������E���t}����x��\6:~~0�b�8i�J�r��~c��ю���p��U�:��Qn}U��^�D�P��mOS"`�$웾�'F���E�4�5r��G� `�B�Ȣ�[;�=��:�[����[s�H\O���Tk��H�Ա�J��/�6dZ��W	{����O/���x