XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k����:����"n�U~Qh�!�M��%�"ء�s4O���"�lI{�һ��Gz��s��P�&�oq���"s����w�u�ƻ�����C4�V� �/�\L��Ľ�ӛS)�tyӾM/{�&
P�檎�#Yկ	y��M���k�2�q�j�GfsW��r.7P/C�!:���uB}�?aDat������Z�?�U)e���9a7<Zr�֍&�u Wb"�#�~dPw]7آ,�םH�y
V�t���8���(�q���MxӔ�B�L�[$т{��)��UOM'䢠���F��|ֳ�b�Q @3�����ZRj6sT�Ò`n��UF��x�L�Zo�˘���4��(�]�[��W�U�OT	u�Ҭ��Pv��k�s.9���A�-�V�a�&_j�ȋ��D����m%�Is�����7d��W=%TM
6�[sd;7����s��v�̎G.��0�a|遥q�(�V.�'����G��/��q�t�ɩ ��P!c��H������Q�>�:�|1#���m�� ���V7���;�>�!��B���`/'I���ץ~ˍ��D�
9F���������r����&h\}Kl�wd�H<5�l��sc�.����a��]o�'�H�9��&3`ؤ ۾�������$�މ���K���X�yxM��=���>TGì���#��Co�=,Z����Rݛcɻj�.9��#�F�I��]��ʩ,��P^	3��{���_KXlxVHYEB    1cf6     790�[.���<RZ)M�����.vЁP�ZV;�1� �s{��O�v��ܥ��$}�3h��S���T)���-��ϥ����r`7�#Ԝ�X$6��$,A|뼖��:L�֪Β������ɋ�}6��5�����U[b=�|u�٦=�m<_M�r�����uˇ�4���j8���!ll�ފ�ي��'?�e�F%}�0�줂d�Ud%��/���ή�t���
O=0R��>�����L/�"F�n��N�ӹ<��1��[se����%�P�PcG�K/����:�+=2rNd���y��:�t�O������
u�zf�<������ԥ���&	��]�b�u>y�-�(_~6U� U��hzƍq��
>�":YU�ur�#����A��P�:��e�x4\�ej�q#g)U�?��W�����&'ύ��+��NS{%l3�����i�g�nk�#�t+jqۛ�C�|���܁�����_�M;l�g���/�Ly�$H�.����{�,rwn!�Mb��PM�<r���~Ҩ�Ƽh�x1�%�,b����GT|��B`���1W!p\^��1����8�ѭN���݃$���	�|�-�bp` ��]G(� ���;��7��zb��U�����lU�P�a��Uւ��*T�	��?�F%oxjؽ0�njH4g�� ��Pa�O�;W	�����;S��W{�8	�[y'������i�f�Ztfm�o/���SJ��[(�)�E�/
�+U�딄���wLe��&�v}�qe8�	����8<VJ}T'x��N*~{8�ɡ~;�_V�Gj����}���ݩ���8�!�7�����[��U4yE�����+�,��-�[��-��:������t�j��16=�I��U���)����D����c��<���>T�Ai&�5)un�^g���b Zs�녍����+���N�*�к�wt>�V�J���=���e���v��&��?�dw��H��V�&ߢ����6�QJE��Õ` ܚ�Wc%rv<�` %�,W<'X�b��3��DkYz�kW���G�Ω@`۞\�y�)��R]>�W8����\��������ۡǿ���ƭ*�#�!���Q��u�=��Vy8�q�S)���%�pVo{S�x�q�� ���Z4E2`�-��m4hR�
N��˴�g�o_���,I=�'����Qn=�fȣ�,=�4���>2?��MX��Oe~K!L��u��w���p/W.���BȘ���idzki�/bi�u��d&c�tsy���X������}�"�*@����m�X �q�c3��Q��d��?].�DהҸg@r�"�������ݤ�)6�O��/:��3����z�l���*���7W҄�I�h������  ��g)-���UYtX������ t`6��Bet�Xz�+���!����r�$��'|����&���ri��{��Y0�3r��W�Rc`A�	�x:�r���rU��M���
?L���5s��'��B��0"F*co�m]M�^�u�-�ý���i�"��"�+0��kMGg��s �<� �mx�Y�G���=ܕe����k�Y�,�����t���_����Ҫf�Ų�FS���gS���f�]��m|��]C0�B۹O8�H>X��o�a�����L.��+�HA�����sçsp4q���%�r�ǀ]���A~�pqɀR�٢���6�������s�̭�P��l����̏�sַtX�d�D�@�]��Z�^̾��*fI�u�.ȭ�������\��it�tYc�:ԏ��!�1�}�&�טFK -�������ye�V�́�8�9G��O�:ܚ�.��Ѣر����-I���������Ji@Z�^~�	�X�!�,�