XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]�%j��&�x�=�][[pR��\���QUG����0�-���k+N6}U8c>�]�w��Aޖ���6�R��נ:r�Z8������"HE�f.\S�	��4� Mng��X��;C&B j���,ս-�&����֐���2ؗW��,���̊沪9�N�b��Ɵs�	��W��)Y�g�J����T�XS �����L6r1���-D�7)�$	��_�?#����<��M�(Q|�1o3Nճ������;��%`�J���OU;y.͍J��5��őw6D�3��i�K}��z�J>���cS�K���CC �F��� 	B�(U@��5� ɳ�g������ ���IP��C�kHؤ^�o���^:(������>���)�wϯG��C��~�dv��xI�vG��L�˸kO٢E7@N��49Z�sc�N�<��w�GMmg5�]g4�xxh���eTU�	���cݑn�*Eݣr��N��h�g!���7��tU4ME�f�-�%�{�==U.��#���g4 ��~{o*e��kT��<A2�
�f�[���V$n�B�Y 2�0
.B�U����0�Ф6�k��V���m����31�m
@����b)7o7��Y.�>�*D5���P��՟��1�S�D�\e��s9��'05p+� ���O D��	�v~e�5�f�c�:�.�"!HU�7ܿ"KEsH�c���M0#���Ү6��,�.����GZT���М�?�4:^#�Ut���XlxVHYEB    1cf7     790�a�C}�R�}a���]�T�%��������C���H���C � A��yT���&|�	XȾ�� *b�D%���h����K�tg���2�bWD�)��&Q�����w�v��V��j)�|t��j�K����R�y�'g��_`��xhk�{�]�M����"����}/���G�J�}�D���,`<�6��r4;��T	좭�z��x'��xw������ˎRU��+�����U "�Ms���f��qp�1���ݎ�i{W�cEB�T\ܮ�_���n׿�nd�p�֦�œ�K�jk��������)��E�"쉩ftD#��L����z+��*�"��������6n��	�y�e��^�#W�Y�ֺx���"�:Y���">y��BC��@����z7'_n@�z��� cUw�UCx�%�tQ�V3CD(����V�l¦��
R���WcW�E�i���g]{�F������=j �[��F)66�_�z�"�0�~V��/Ԯٶ߂�;<'t&�`�ӯ���<,�&u,I��&�%��X������.�ే ��GF���Q��iw�x�gQ"ʲ@��P�18XV���qZ�?�)JO�0_r�|@/��hc�;��^�L�6Ӑ/myik�����0ee�a\���aZ*lG]=���Ρ)�|�X�&�*�]�)�|�����/[px�6�e�uPz'��0rǉw��Ic������á�E1l�L��D����P��^8�Һq8lJ��)�3��!���u|�P�e<m�]�bN�:$�+���2B���$}���	�z������� �ģ����t����έ׽���sPH|�D���JBC�r��zs�S��v�3�;�����
�x�,f���s�������an���=�kU�	mK���dd�8y�xu��&������q��R���.��ѫ߀�̐�ƥ�����`��n28�V�:L2XV�&LRA��H
��|K�c[vx�stu<�u�Z��V��T^7��5"p�қ&I�W��]���	]�����)��G�=!� ��,�=I���"�r�5!��������v������(��qe��xm�~k�Д�;Wh��2�r$�<��VՁ��{R�g��2�Ƚ�����%@�_��G�=n�`(�?�^�f�d�)eb��p��K�"Pp*17��䧋�Om=��zF�!Z�r-%�T�!EM	����δ�t�	��".>�,=MF���4� ������쫨(�]R�M둬4�Ew����M`�����z�|5uV�t����J�}�LG���IZ�s��$�[l�3e�k[^�˿�!�?P��%)�kO/����)[ط~���R�vhо�̂XFoPe?8��3������A�|'�I��6���5A�B6� Tȴ�������E���[L�(���,���;I���O|kg?� LcyjI�Aq+�DV�-�:��b9�jg�j>���48C�!��<d�)W���F����*Dؾ� E��U15���V�>`F�P�s4�&��Bי�ar^�z��`���P'J����f�N�5���G��J@f�����R�^��d�
a�y}ع����Zo_6����a���3����7���x���E�D1�y���yt�{Z�x�/���^�Si�BW|�TɃ͌B��Ă�Cu���ɕ2G�� ��'�в~�)� ���f'j��{�g�T��X��ࢵ�c�<[j�~
��媩��hۜ�J�8��cC;�d����W��*�>��PX�@3Qn��>  E�w?�x�����a�3��0�c�I/i����U�Hk�J6��4���_�$?��sIY�h�sp*b�,������â�P{��G2�