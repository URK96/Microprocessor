XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���f[ٕ���b����.3��^�drA-��(��5�Y>��F0u^j:'G�Ax4�[M!G��#����\(��z�!n03~,���W�ضa>�!�z���<��q������u=���Z��ջ/�輯	j�q�d�k �F.7Z�&�!��Ɉ�u1��$��e�|��� yQ��	6�����ש�LN���}����~���5�eN��LĤ��9A����I�����ȮA����ɬ/�M� ��VST��7��GG�(�{�����vux�c�M����v��Tj�9 v�
b4��������S�}ڕ�%;"ci���`1p�kr����~�Cc��8:%����#�A����'���^�5l|�+:X���.�a�*��V�#��X�t.n̿�xL6�t@���u@�鞜n����B!��má���tS+"�6�'
�ۍ��9��O��#��06G���x����'�����5G[��L�w'P~ܴט}����m0���0��/��NqCث2�>>���fB���1��ƑpgjجNVV>�p��G��W�3 A��<�6��wg�+�er����xuP�D��(5�1���
���?
��M�?�U]�^��3+�r>�Вj.�*��T�yl%�ˋ�P�	*��x����i���8���9�a@)2���Y�,��w����m�*�ѝ����D��C��px������E�_o`O�rZ[�@H��'�D��Q&h��U���XlxVHYEB     748     310��r(f�F�-�S]�xܩ�~#Vr�yL-f�~�I���9e�Δ:DBQ��Ē�V��R\��C��P�\Oְ�gҵ�WlÎ��w���͑�`�XX��P4�]N��N�� R��Na>^�2>D��:o����F�>b��CW��Xߍb�v�C4PWV��5p�TKm�>E��` %���n���-9r�������2ާ[|�=2�F%��]	^��偡�Դ$7f'm�FN/}�>eJ�� $#r��y}N�`/��p�x���{dd�&h�Q��V��Wl[�����LGE/�(��\˦_I�tAnZK�".x��W��χ�1m !@\�8�w�ԅˠ��1����H��i5��?�S�*�a��(��Bn��p��n�M��Bsn��� L�q۩w�x�Ag�am?�/�|����l�����D��V�wåZ[��O���F�Tд0��6|��գ���3g>H5 }l�7hPCh�&�YJ��oW��Y����	ZJ�6'�����#���^,�������4pB�«1]�5vM���'x�yYɧ��W�z�+�����EQGtW�4(M�^�tJ�n\֣;�?�d�I�PRlT�&�w�C�C�΁K=��PA������� �-�C>,d�������L&��k�½�Ş����>��Q�ct乼�|D�k��M�Ãpg��k��Owك��e�`������W����7m����Pb'��ٲ֍pT"cƿ�� ��9R�J�I�.����X��w����:s �*