XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���:���<�r"nr��D���j�,��y�H�7���������G�����y��5�a��Y���'�t�)u>������\��BR����yY �n�h��5Q��#�3h;�$�g>$��l"-�r�rIP��3���[}�I�~ )Ey 3��r�[uqC�B�!C4G��P�U��S��'ԁ��^`�)�˚����
>���@Q������~����~��L,*(����� ZN�.�8�#����/����7�w��Y�8�3���흥D%�Q��s~���;ޭ z��I�_�,�.	ؒJ�/^S�:���A��y�q����k���^tb{	0�;���k�d|��X;����#'�U"��Jq�1����9�I-���4�Tcš'�a&ʳ�'�@)zU��詴}���dl'q�0�����!�>�޺� �������-()�<�z�q��'ڝ#Ͱkͳ��t�O����?|E���o1+�r�O=����=�lc��~��+چS�������t����h�����hy��F�B0�
ZX�;�D+���يT��d�0}9�����D#�"PHB����}+�Ӹ�� �@�e$O�tno<�a���k��?�!�����s$I&P|�-�^�Y3��vT�XD�w��4җm7�-��}o ���5a�왖5�<�D�݈/G�U�1�:Y��y�v�Nl3B0�A����a'�Jn'� «{�A�@Q��P؆/Z��f�K?��f�J���/XlxVHYEB    1047     4a0n�!�@'(%3VO�S���A*ܹ2��dE�PjE � �D�P�ku��^ҭ"���ҡ幭ͦ-�p4�_��eE�h���T����޿&�QR�E� ΍��B�1,'�rܞ�{_���E
�"D����w%	�[$��c��KtW���Oun�ޫx%��}�3�9U�Zԅ��5�k��V1A���zU"�^Y�;aҵ�ٚ{���k��z��*Ƹ�5�W,Є��4��q,�B�X7�ߖH&)Gih���-!�ͤ��
N#�B;���`����"���^r���P𔝄$ĥ}.��+���XFA3��W�#HF�y`��e5�3-� W&�&{7&�FV[��	�	��V�vW�}Os�� ���L��@`	�x��̴��.d�S�$�$����1����8����� �+�9Ny�+�2�����o�Yd�qE䯼=��̆��~
E��P!�&L©߽��-��"b�X��M�%�u�U��� σ江���ܵxJw�U�͞H�q�;!
�T5X��K��}X��r�8�7���qs�?Hl��~�9 L��f�|zD��D)i�A�S�Zi�FC���'J^��v��\����+�����['�2㧈�����P�'�ofyׁ�/EtN:x��v@qd[����R�9��v�o�B%u�ֻ��y=^��w��.�`�H8�"OH��Y���bX������ �(���,�Yq�=����ս�a����+t1�� �����"s�>�y��r[�ao�{���z#i�<�'���|d�j]�\�4�E�x�C�)�#�	;l�BkI1>��9^��,�^U:\c���?z�2�)*v�+�E�6�-S
V n�I���g���~��(8E�A+T�u��u8{�����N�i^�ЪWm��Uz»eY��r@�k��Is�9g���Ӯ�>,�c�F.��hsF�d_7t��@9#!}%�`C6�^v�r�,����s����.�f�����N�=ݻ�6l8�%r��6�ݞ޵�O�3R����w�J%THٵ���	�7`GMUb^@n �8�~n�Fj��x)Ď�L��b0]"�V�5�FԒ�o�o�����˙�yn�Re�?ht���Z���S���E��&�\�ޙ&�i5��g"�֏XD�3O��|,P�҄>� _�v��3