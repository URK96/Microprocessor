XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����]T�X	l�aE��M:qU���`=�N5
�Doq! �]�@F��!Xi ��% �W�Wv��1�6r���.@� �,s�� B��`Ot�Y����S!�mRN2K�3���rF8q���g��~8*�=�`�׎���+�?��5�M�g�o����RiACu�+h��|Ye�H�G+*���F��c�A�O�j�����$��6 ����!������C�4?[��6����F��Ah2�.qNU�0N�V�R�����_V�/l�k�~{�������&�j�U�a 6$i��ʎ�[���H�Z�N��y��?��?���ݞj��L���ĘLps�3~����)�O����%�وG��G�Ϩ�ԍ.LZy����О���-o^;�I��w�<5#�{�~�o��}m��6~�M���7҈�_�2��O�
�=c�
,�b���k��8��xݜ�GNl0~0�~�Ԩ���2�W;=��ʽzɼU{���S�*�x�bm���H�Un�Y����5�+�qF��<]/YոA���?���F�y��M�	��WI��MT��$z-��JI�pjg�����Bt@W1�~�nSGh�uV9��Ra�>\��}v���g����r3B���G�K��쩨Bx�"�n#ގ��k�K�O��X2����R�S�`�V=�UB��9�v��@T��ٍ2�<�w��3s�sD�u�Eb�*��;�L�Hf�0o0}E��)՚�ƞ��6�ä�x�]X��u7�W�e���!�9bҬ��XlxVHYEB    5ff4    1040x>���y�Ȁ��08�V��4���=5�ω�y� 6�;F�b|�}��0�� ڔ=�*��J�Z���LI����hO�Kh�z�_�1Tu�V�pD��T
lmD����r>�5r��ȋ���ĭ�e�� �l��o�п[�G��_�@a>�s���(4dnK.ۋq m�h)Zv����߇��1b�C���Ę��d��^
~c��n����q�Iu��܍�-�hVyx6���-���� �6��R`M6����L�pe�JT�F���*?iGe=	wSd�H.��l�]�ו�b}4������,���@���-��SPY�%�fEkO8�z�|մ�԰�!�2J����Zi��;�o�r�CTK��6*ğ���L�eiȝ4�q�d#懁�	����Ǫ���/���0; o�W��UT�.�� �EC�� �T�u`͛���V��|���Bϰ¬�F����
G���֊�A�
�&����W�~�l^b^)�>Y6�z)p�W����A�.,��F�F�3�(�H�,=H�h�3�	nqz��@�����:'Z�������VQ�ή�#��*e�j��u�}�]\\��.6p�~,B���A6X<(3�]`0�$�C�q�v�k����;5�a�`�"h���C��[��'-Q��]�{���들Xq�m������W�FV�x�%LT�7��r�W�Sl��u�2`��S�����@��TDjj�u7;�m����@�w�[A��O�/�q����������Gg����G��gy�b�8���z���nC/�9��Q^`a�-�!D�A��Q���ƹX�P8Sÿ��6g��@���|�f࢐P6`�mRj���ڃ0�p�c�)��OVj/���t��9�O	\ϭ�x�Oۈ��/�A�	�d*�]t�>���DGC�.�6L7����܎��?���}J��?�� ���]Q���tk���l�G�f)ts�B�A�+*k<X��a�Ù�1~g3M�,�p��c�
�Ői�˃o�<��5��8�jY�:��s%�0/[�Y�@B蕷u#��s�0@���Ir��5 ԏA�H�\�N@5/ݗkTEk�ø=�A�N�����'�z��rH%���];�W�����)";r��x{���X>E6����;|"B�"\��/�㫳w��c��1Q���8�jX�S��@���e�#�_�!h��}���ε�*�c�s�:���v�Q7��P%$X2'�\����ϵSg0ʪ�9�R;Eℑ6�q���<}���[�7��M��ާ��)��>�y��
K�ӣ�&s��x*V����2����2����\ 8<��o�ϩG����Ô����Q��+�-����.���R�#�b��Q�pm�{��?���y���:����k�a�\݄��o銀K���q ���~��Ӡc�'y�S�,tQ�O��Z±	Zy��y�ێ?0��\X+�Ң���-�('�ٓC��AX��a�:��m#��@-b����4�F��Y'�ڝ,�;���'���_U���BQ�P�G.LOM=�r�>��N!M&Q�C[���"M�(­jO)_l�@`z9�%l�nt��J�H5>Ari^�dq~��k��w�ә��!Л�
��=��޽' 0�F�0���W���&���Y(x'�+��[�R򋘘�o�M��$��W�V��@ŊIh~>����B��8D[}j!,|���`珑�C����X��?��T�!#�X��	�F��+������
0�uI,���,��1�=H)U[�!)H�˖�~�;�y{ۇ�g�����u���ܷ����-m+��o�������������JF@OX�l5�<Z�z�@��y���ɸ�bՂ���w+���oP�"_P	G����;�;��l��d=5��Q�?ia /���^M��S���p�8K�D�5:Y`%��z8a��4������0;)�J:�Q���}K��yB=?�Ĳ��7,��R�#P��3(��kCƀ���G���S���+�ո��|m����3=�� �U�)�٠���!�e�r��P��$7�\�c�~3;�G�+�y�0��O��2�������Zó���u��vv����R�k'���x�r_Zy�z��/X2�;�3Ʈ��Z4F(���������В��v�Osõ�����0�LM��ldU�q���B�'?�X4q�1��,�)� �+dl��-^���^��N��}�����ƛ��Y�H{�$V8sݡ	;��޺_޿\
"n�쵅F��)Tss̺���$N𚣔�@������>~�xm�j�ez��6O�z�C�
Ϟ��AݍEX&�O���ay����/fR�CؠTR��k�G3�&�Tø�3���SQ���f��46-" izB�
1LY�jr��l�ɯv�p�\����Z1H�Gj�A�~U�O� 
 �`iU����%z���-�O�\�7h��d]�T�<}��t.}я ��ʼ����L<���sB��c�U��٧�;V�{�lg��7�È��ѻGd,z�A�?�*s0 �2ŭQ��xr��<��a�ӉH� ��*-9�ۙ���(�:ꊄ��6e��v�$����󡳉=��o+ug��q��Y>��K�0��(>�/5�0V���$�I��==�SV��pNaq
����g�_��W�0�g/��6�9K��/=�16k!0�W�ҭx��!�Р�M!@����r�T�r0�!=����86}ץ�tB˗i��X�m�����Xz��H�b��C��e�dHR�zF`Bc�&x��N`�#���g`ؔ�F+MToz_��m ����e��J��v.���d���g^ʊ����3m'�&y�'.�U�gBA����(�Q�EcKvo$R��w���VQ�{�2C={��V��J6�r̫��Xm��	Q��e�����!18��n��I��[�2ft�_tL/G�c���R5
�(����u^9}���U�&����R	�c�1b.���#��eX�����F�6>�,�,��7����N�ۋX�\&^`j��!b<��� l��bN��F	����� ��-n���@�8��:��]�rY�ͺ�����e��(%����~v�l�v0�;�:)�$ 0p�{� �����:�Y�ۈ�II��	�{�V�Qb��K�98Y�X<��2v'���@��?�������#i&���O"tu�d�#"�|�^1L3{s#G���
��F�P�ڑA��H��A;����+k�����>9pF�\�ȮWTl �6�𢣉L7����M�7�(!��)'�^�O������}|$���2a.ݨ�9쨳l��}"��3���Y��̑vR�>4lT[²*s�d���+��"0�t%����#��Wt����oݢ�0W�:��q�4g�6�[&�j0S�b����I]�[m0�V�U?y�����$�,<�8kr� ��&�S]��E��}va�d}T	¶�ķ0����*��<�ԇs���
����:���$�
���~q������yq�.E���lړ<�*��O)�_���t�_�A|b���6K���mf,���K@���M�mL���2�@������	L�9�(��jQƸL�O1:I�<��|�������s��
�$Ԝ�m�J �*�	��FC��Jmy1��u�yi(�.mdS`i���!}��v�6�@Y�(�}�� �׃;�}���by2�>�5(��:2�C@�Ɗ:��F��JG��A�U'�}�����H����ά�!��ݱ2�`Z"[v�!���q��G��&I�Ji:�yW�U*�!�;��D�Y�cg��� �LcV��U��;��"7f#w>;��'��U)7Ν�{(�v��b�b�F�K��+C�x"�_�4ƈ��_X�'\5���tV!�%R~�����w{�{Z������/�X�Hb~Je��^�	��Œ�4	2q�Ib��B�<�+��6f� "�j�{Ğ��_�@���z۰m�U^2�^�e*.�y�*n�@7Q�x����������;S�4��e*k_�؋F�s1
���Խ�Qo�*}L��2Q�&���{��ϚХ���6��ruQ��B��