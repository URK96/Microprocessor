XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A#N�uG����(�5�����ED;T�Bf�5���8Ȇ��Lp���)�dY�3�U:��:rF���w����U�Y�8ǐ4Ǚ�^,����G�4���*>�ʖ$SK�n/��8].p!o�W�pX��0n��g�d���9�T3���-�M9!5�[����Bbh���ҙ_��C?��:�/JH�ʧ�v���<ڤ�J����|E
��o���O� ����G5b#�v���0�E��߱y�^O����v	�x�cJn��� �(�U��M}.�I�,M�b�ƹ�|�![����e��JW�urq���S�n��e�K�X��$��薳�OJH/[��u�u� ��N3�sd{Ұh�tn;ߜ!`��U���{ K�����,��Ƶ /�p�o D�F���B'K*�d�)r���S�{��/F*��Kf$ӹ
��{2,?�$�f�/��0'��߯�c\�l��$��%2��W�dѼ���M���;S��@��p��e$�}����8D��I��F8.ag%����'��98$�s�8��u^~��Hm�w�/����
�ޅ�+�qX"\�Du�T�+����J�����i��W,�J�~>��2��P:멛#l��Y:�4(��󥰃øU��M�{^����[�(z�����4���л�?]����8y��I�����|�oF�8��Y/{tt��tC<��
�f_'����Tu	2E��x�hfI�θ�|���K�R�\���J�$R���7�'��� rv���XlxVHYEB    4a98     e80tL��̫�FYo^����2N����UkO���ó�1��<�&?/��ڣ������9@v$58���F�<.%�%��F?�Ԁk!�j�'#��,�9�#����S ��Î���ٞ�N|7�:����)��j�� ��n��b��2±�0f#�DA(�X&YB�H����O�mƵ��>��X/�Y!!�*���C��p�|8���ze�͂��G��^�0;�h������i���#�B�SB��}x��q�G�N]���B��΃䓱4c�/@��P�7��.)Y̐�f[!靕Q��酼��Z�NL����\��}�K>|d�X��u��.�C�I�
���=�V���H��K�}���s�jG�G�j�D�U�/��ҫ=:��`0%�x����Xd�ްJ����J�;�k^����(�7��Ԅ�̠jR���[���Iމ��!���N�Զ�Tl�"w�� PY����$!W�>v�H�ϝ�,
���H�5_P!�D�6L��$�����W�+���v}YH���4�y�Z����Яh��Zv�H���d�Nj��p�c��$#wHE$�#,Є��E�Z�퉵ۈ�E����.����.yG*�s�+�)l��%��]5��T,h�� ��|���p"v%3�UX�+u�{�)�DT`�-�Hʝ�41�x�`L_���ftޞY3�s��;� � �V^��mve����@����~Dyo7�v�=]���q�'ᖕ�m�1����������?�F?������ڟJ�|0"eE�)��拇���6�DI>+!��V��8'�γt[b��A��;)�h�"�S�Kطz{��O!���"V��J��hbVچ7�$!j��wp(�6y =B/�@`�xO��U�IU�`����o*��t[
�@�no��D�s�/�=����c63�|�;ᇕ�u��=Ro��_���yRkL<q�ѢL�4Q���)�0X��U�?3DƖ�c�KIG�XB{{���>:(v��vk�Q�qq[��ڙ��r0s��)���hꇮAii��粸��
	sK>}y��=���ڵ:q�!�����ϳŸ�˵JAJc�I+R��W�d����[s������$��@�Jf������f'F*?��kGi/Ze��J@�3r%���5P���do
�kO��^,ި�}��Z\����͏�*$6��+��	�F�#�����ꃷ|��8�U	_跠L���Ʈ�f��-O%3x��j��-��m���QC^��ӑN4r�>"�e�,����4w�Mh��YՇsU�;YL�\���Lg�τ��h����f�� �����[$�Eόb]��Z�E3�y��&V�z�g���@Z��F�(	L(oM!��n*�^�EM� ȶ���`�/����{1�+�G��+n���AXˎ���`c*���? �4펮0�n�p�QwBN��6�%M�{�؟�+�K����Ϻ���y��@"CH�R"H쑌hJ��r�z��aL��L>X ���U������b�`j#�ρ`$U]�O�b�e�t�8gKd�]�I�.�9gm�zK�h� �(�
�j�cs�{[AL"�N�i�\�A��� @:��ؼj3�bvw�@����#���H�/�Ufx%��yR��m�r;�h��ex�TGs!'(}��+�vݔ����6/��B�s�	=h��R�ָ
�ds��y��9�t��h�!�"�����<��	6�荸����%�n�E����djp��`F^�X��h��!jU�c�=!�N�����f*�Ǘ��ӵ��(lol�ǋ<����D�$�%WW����`��#�g�x���y��=������4U[~�lc�bڱ`�"��V�|9�����S�C�ô��y�bEX"%��,X�!P�6��6��q3Hm"���)����rK
��E_�C��7`�bgP ��%�ԏ���= 7�5��Z�2��>ЧHj�5��O�|����E������m��=F#BtY2L՞��&֦��j�eԱ��[�i<C=�vB
��"�$�@�Vײ�Ȃ ���-�Np����z_���b	Ы� �%�v��p��I¹陲M�6�F��v���_	_����c��{4�~�N��tvR[_�	�p���(���.d���{Dq,H����\�(�m�����-.�
%}��s�-���3�de��?o�����{���`a�V�[��AS�--��	���X� K%��D�����v��3D����@B�+���_/��Ä���zJE�$�{S|������.�9]���,��Jl�
?��i2tXS9~ S�fǱq(n��Qj�+n4�+/�R�&��&1�7u��5?�[ŵ���h�ٖ��z*c��َ瘀�q�GIY��gV7D(��]:���2�咝�m��lhW���94ED@��*]�	hT�*��`���!�p�'ɒ��%�-#y�H�Ŀ#a��E:.��MF�*3V�i��v4�����uG5�'L��d"1�Zt���Xy��W���C���;��C;���fح�L�`���f��WR�V�p��ܤ�A���y��fv�zj}F�+"?�Iʘt����2uWU8��gͦM����N`P/�T�\T�L���\4r������O�o� ɛ=�^햑��5�ٱ��k+W��w/h�Q��e�[Eu�����^�}�l���ؤ�����z�IX)��nc�)7�5�B�2�ދ�-ש]��7	e�*F\�.�,�)�x��ċ��κрF�M[��)5��'\�D�،��`#\���es8�۟(
���o�U��0��jH���I�C�S�yQ*�a���Y��ԟZ���B�H�c�	'Ӡ��)��2��E��o��p"^GC#R��}�
}��:�����o���^u��/���t��J���+�0�!{;����'��hN's`���U0�����vu�7���
�AX�TON ���\��A�bAi%+mV��zK�A����&b�_O,�ڨx�����x�*;[ԥ�F�gH��2`�d��)��2^x<`��D��
��ڜf��-�u"��(V��g�9��68?��Eo�	��Y�(�U^c�ե~�����W©�6�[��syΣ�S�����>uE�����{��4���gSAOg|+#N.�� A���X	r�t=ܘv�V��mjCKE��@�0I#8`��y�,M/�uÎ~�uu��������ch�}��t/(�s��w�7����!��ca
%>��g��Q�d�7͇]p�<%�@�-:��j�:D'��yB/��um�z����Px�ޙ��M���h#���K7�oE;��3��gL�o�rr_�r}tV.:6g���]�%�rv���/���9�M�$�w4h�������̡=���q�8o�H�7�cYZ�,o
h�Ȫ[�D��0q2����Zsc�J�<�2|��h�?x�0�>y����z-�&�,�S�~�Ҕ>3���4:������P)���)	)����ͪ�������G�����]�X�ϔ�	EJ�i2�P�*������T ��;d��0ca�VՑ��F�k3�{A�o��*�g7������>h�p��Oq�i"���U���s�="�