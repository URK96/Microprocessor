XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_��.l��݀o���RX�4���)�Ir7����
���-F��Q�Be��Fg4к6�ژ
�R�����$�q��C�ʦlGg�"}��V04��	�3Sű4�8L�,T�h����Ag ��Cd�(���j(����Q���%�1s)�Q8F�ʿk��Iጤg	e�ډ���2�@�"#�-K��et��T�A�σ<@]���r��S�5ikd3�X��~Ω�E����oE�ŘB���=�J��6�i��g�9��[�P�V4��)9���"Jv��eM!�#<x7��|�#C/*��;l��5l�n��d��m߷ݺϨ���mG ���V��"�Q�������꽠8��v�|]RxF��!�EJ���"�*4s������Q��G�<g'�Rᅗ��O�2���JA��U��݌�v+�L{[��O7J^�/m�ydff�o�q����mBc�����0h�LR�ɉ��mj��ԇ�b�ø☗�\�
!�Vo�AMϒ�=�Wd^d��c���Y�l��usZ�C�ymԯL�i�&.���ɾ��R��-���*�?�]L�G�~�'bG[�t��4�$�������(�����%���]r_�(\Vz^;5�9��+�����j�,l�:�0��QRs��<;�^�a{�]9҇r�(qo��¸K��ނ���5IZ��*��\$���^,�.�j�ˢL�W�������=M+zI4���d/��7(��?�"�L����x$8G	�[/)N.}IS~:IXlxVHYEB    50aa     790'�W�s7���e@&j�үH)��2��3va��X'}x���)R��D�=��R��OA�j.l�
*)��L\��D��i��=?w�|\��;�[�@N����4�����s��V�aF�cC���|�_&6�N�����Qc)��ů*��n !a��wR���o�H����$��ϥ#}�)tp;���銜�F�U�b�����(����t�ؐ0�N�d�%�cG��#DBAd�̊ٔ���*�e�r��{N��&��⯫M:LxrIlx��vA�����b���M���~�z�ů�\�"2l�M��f�c6\��!��X_z��vn�jt��@�Hݍ-�xT��-����������l��lXF�U�E���=��i_m�1��ʅ��o�N̏����V�]���S�w1(�����/HLby�(�]�
��G1!k�AF�bMlz�`�r��Z��*�>D�_�v�,n$h��ZϜ���< �,�Z1�ga ������P_vi��Uo}Ҹ
�Q�QJKXD��1� ��?�<�9���谱K�=��d\m�o��l�X����e�+��cw��F��dS��Cs�J��y��:i���۱�8����if�Ff�"�m/FVC�]F%��t	,�w�� ew��`Ӆ��z|f:�����X�����(�q}ە�z�P��Y�>b��n�\���/F:���a̲_�Ě�N����P8� Ոy�B�4I����[|��'����;�5��"H�(�Ms$P�oq-x%3(����ϼ9ֈP#�Uh����K�J�=���d�aO��6��k�d8�7�	��W}I߇����5�mAu��؝���#�q+5�S���?Ks9�*��\��� ]0�yuy����5�1 DK�K<@���:�nbo��)|q��deM2/�:Q��XƱn��(��`��3�ġ � F�ed��Y]O�|��u�y�s�����4�QO.�T�u%nf�!q5�����ͅ\�NPP��D�4_�ƻ2��vlJ�)-xo�ދ��� �.ċ�"
�].;+����	�Z���./\H�$�E)�*�TFR
p��gx��'Dl�慏�n ��T_iӌ�&�2QKv)(p`c.�����
#c3�"�W���%��g��@�1.@W>7��DZ����]Tɼ�AT7����bGݹb��b9>.�I�iPڧH�31�B�ok6S89gĊ��L'_/,���@-gB'�ܛYZ1�� ��>p���l
�"KUj�2YS�8�GD4,��]w�c�|J�$z
�0,�E!��0�j���ɧ'���dQ.��?��X�c��^c'�]��8%�� �/>�M..�
[��}^d���@�!�Y�
"լvH����?���Umf��#"p��A��
]��qqLg�!?M��38��l��-����S�ɴ�p��s�ٗ��Su��k>�
ߛ@T���Aw�0qjTO}�5$�E���J�����owH�ЁBCc��Vչ!-����YbP �̏�**�j����[��O�`nܿ�0���/�)�~�����"}�;%��=�+������&��n`��G
�w�#��D/���Y���W�,̓�ԥ��������O+�b�c�ZeC������p���`�Xz�'ԭy^k��n\H�T�I��8L��C#  �R�F�H��^ؓ�D�Jtָc�hQNu���\g���X%3Ӎ���
�
��� *9;]�e7�kR=�=ӯR�Q0�ҡ@cI����} �-�:��4bҤ*f�>@�Q:_�X�J���aF��V�>�%�|/��ˀ+Q����D�(g��Z�(r�E�2�0�X�/I�6߄�t���'� ���o��H\ã��WzVwv��u��|w�i�kRg2i&r�� ��R��l�_���l�Xa��;5�
��a�