XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��vLR�O��e$�$��- �{Y1�����r�N>��7T���>����лMl�~R2l2'N*M]��h�lk',ˠ�Cx��!��&ï�įg�m�g����e�Ryā�tA+����>,8;��5|�*�Q �Ű.|��O���!�{z	뾽7��<��7}T�<�:���5w��z/DM��ht����7�&=Φѵb׆��*��K�B�����8[Q0#g�bV����͋]J�e1��µ�Ǭ�T�8ͤ��D7�F�9��U%	 �G�/R��r%���('��kTW�}h��|-ι-�t�s�t��9���O��|�sK�2�'��ʻ�$	U��vv�C�<�d?F^��E�>ktй�8^���o��Q�N�k���`����.�7N�K��t�
)�g��2Pȗq��M�yW�
�i78���}��/����T�qyQ�I�� 2?.φ"�E�r<p�ؿj��dX��c���CÝ�t��~@uJE�!�sۙ5���� ��9�h��4���� �汲�7h���8�e��eV�qY��Ň�+�2����|vj��1��cƪjk=v{���wP���H�cFT��}b�|��H�>���QbO�B��t:���D��-�Ԃdv>ĕt�_w�N�2M�G��7��Fh��=�(�4�k�.6N�L�2�h݂�x�����a��n
�.��Iۉ���0s|jgI�1y�D���x��Sop�2�y�"R�\$w,�Wl�ǎ�+9코E�32�XlxVHYEB     730     2e0�M�oǞ��`sz�K�2>�x�:�)�(ըdx�D����G��bo�ESUk��*h\�
 V�e����^�]���<h�_��`�Nq�{�9��W��b�L�ײ��N��x|2j�����rr+XF�"��Ѡ�����-�$,w-� ��D�=��iXZ�C���� V�}[R�[��f��spQ�!2�
=��x�#G�2�'O_ÊP�����j��.X��"��N0��U���;d�Ad.-<g��:.>�8]��З=�Z��5��=X���W�0�/O0L,lC~T\��-t*C��S�0^����nlO#V�V�R
8*�7�y���y��=�-��hrsڋ�s2��D�\��	��B�o^�Ӣ]jq"�������L��n��Hp�V� q�5���>��*'v�����y����J(�%RjV�����r!R�LO�gY�Џ�/!��7���{�]"
���8�M�w#ȑ+�?��fֈ���/�(����s�b�_i��$������w!�jۂj Y~�ט��#$����T��@�9-۬������G;ʼrЂ �*Cx;�Vd,Z��ͳ���ӫ�Z�"Ќr�f��Լ��{�B���6����p�,��� W���bw1н�~J��ۓ���R�2��ƣ��0�%��rE�3��z~>L �����ҵ�#�-j�F�ZU��W<��oWӄ�c�J�s��-LYb����M<|��@�£���}