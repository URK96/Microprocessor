XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z���Vy��h��Z���:�A�_��ZRu�ۥi.E�mP��p,<w$�W�Wa`ã��e�&��w�Rx�?W�B(q�������`��c��19���U�KѲ���r�zR��C�9Z�~;�Q��*���pK��=�S�'�^�v5�QM�ge��Y����`M�As��o> ����jG�(l����vQ��T����t�]�a fQ�qT��IǛ��fj�ԅ�`Z;7���i�����+�2ң���Ѕ2��nr��㑰z�ߩ]��E3w����u9� H�4x����4l5��u�� wˊ~���P6�M�ا�)$3��8�Ϊ]������6�(]��f6�wx}H2O���(����<r�A�<%@��f���2��or(�)&`�}���sT��g4n�������d�pЃ���Mۍfٹ�-�2�o3�]�GjP��ix���1�a����&��;��l�,����h��u懁Q	�}@�>�SH �1΃�7����I�.[�H�t��D��2�W<�S-=
�rT����"wJg�h4>"�p{��O��B}k�W�/�6�;R�+>m�`�Ԇ����� ��S����)���Uc7ݔ�9ZY��Y%M�����=���q��߯���BZa�y5��(j�D�!2;c/g��.Q�Mٝ���
˫W1�EvJ��˪* NwřLD�x-7D��`DW������QA1���3��bOu����VA�D
r�FPRoL��	�U�'k�T�XlxVHYEB    2fb6     690���h�WVi�l.�/�]cO�`�&|BGL�����0"�y��~��H�m����J�i���U����V�$�x`,�L:�*�{�RN�l�1����ho�>}�6���S���4.Rl�?�>�,�W��2���2Н�R��S%"8�n�Uh�R�2���pM-�+�[��;�e=��9c8PJ�,p� �Q�����n��V,��d���͘q2JG�C<"�� ҋB�!��2qgQ�ڨ��ҝ�-2��`�î|���U����J7 ��Y�Nޓ]�M�V�mvĺ��಻��>��Bu�?�%2����0o$�Y*�&�a,W�'���"6�D���$Q#=�$a�_�Dc�(:mFֺ�x���㤕/:rj3�3��M����H�"B	�L��
��X�f���m+�?��S"U�>e-}���z�p�"���1���4��N���k�EA�f����(�M��G��T@FA��i/Kx�"���ʞ�X�t'dMj�s���{�>�-!�-����a6��C;���*�/7���P0f(	'��F��eĆ��I�\�^r�ZA��)~2�M�@G�3	�1t1*Kr�A_I�U���S��^�?�ƃ�<9.閬|޽�D5f��k�jV�����	�����..t�H&)N���=��B(/$0�a����i��J��a�6��}
�\~l�)����˧>�4~���i��2V˱��R�J�Y�k��e��P2M1�	�c@FD~�,k��r14_-��1D�j���a��0��̙�w�:R�&Z�$aWY�н��2
���Q "�Ƭݝ�>m�`��md�d��8��A��-1	�������*�L��g��Ĺв�ܣ�l*oM%1�-�����
XB���-K���\Z�yg�g ���]~��`ǽP�*�O10K3&�KLr���ƻJ��xf�0�t&�1
JDR�I�=b����7_�X<e�R�@@}%F�����,�e�?�9� �B�7
1��I<%���U{����G�oe���l����_�`�x��JS���sgI�,m=��8�!%�ȇTl�!}.�tT�a�Q�zȕ죀����Jb&���gl�:S	���/�kO8t9q�����ڋU*��H�&��}ou� t�h´�@KA�r�3���#�7�@T���E�D;>�{��?�"'���}*�����I���s~��7P�� ^�IϿq�T�_t�=ߡ�g���� ��(��!����m�c2X���	B:%��
���&�\�Ӗ���yD���#,�>�f�{yF(��Y���
?��շ��O��'���^����2��?@w����-qC?��ӹת~�xM�;H������h"�R���
��;�����r��^���L�>4�p�ȍ6M��򝤡C�"�1��e��0��r|w�#��2�
�ٛd!�^ۣ�|tI<�ݐGZj�RE�[��*#��PC@@_̀Ȕ<Gyʘ��|iHਊ&�?%]�5,	�����],�,�<���U�*�&�]ފ�0E�JE�Qi-�
tQj����Z�*�a����
f��HJ�|�70�{�f�kN}@2{"��1����%`=ݫ������� A#�`4��w2����1�X7qc�fҺ���gg�3��j�