XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j��&d�:`�.����9{Z�"�ع�nH@��.��q���_�`>���2���z���Ѯ��̔����5>����+���SÄE��*�$*����:��aneN��r|Q��)%|㳫� ���;Z�l�G�?�\��t�,�E����'�cm�ߥ�o�����1z	2B �ID3�xM���ǔ����yv�"�bL�1��;�7@�7	��Lc{K0-gk��v)���r���S��@/�A�)�agԮ�����I(���"�lSH�<Ȫ�����0�R��6����w�瑲��ZP]i"�ɽ_p�p�ĵ��ƃ���c�.^˂b�����^;������U)���d�q[(�W�G��M�zcI�"N�,��5UÀR;I;�����9�|Ȑ]�(�Ϯ*�z]Ѓ��4{������>lkF�`��DjŏLkM�L�_�����*]�M�U'~SN+[(aCl4:���d�� (����%��`Y;�����n.����	rd�=)��}���[-'>��.�g��ԅ�eS��zn��g��0&	���{�ԑ�g3+v�a����z_���͹@�3����&�F�6Ų���'kL��q�;M��Ŋ2S#�ՎUV�I��&ĝ��v��-n�R��o�n��r,W���u�a�
U�n2�d/� �1��A/5�{�@�D�P�em�]���~l�~�[e��g�^������������XlxVHYEB    1041     4a0���G���*�M�ğ��S�����G��\�m3��?'��z���� �h�MR�ضd���ô�>B�P�pf_y�a�+���l\�y��n܉��a���J�, Sa`��&71�W��v�+�}ܬ�q��?�A���V�^�����P��-�uZA቎ݻL���P
L�qyh�1\�Q o�XQ<{���l���W?!m&=�wWŅ�1.�����\�)G�sX�q�6� j؃"��#�m��b���k}/i~�:F�z�1�f�'S�������P���%JȖ�Ԭ1���~3����U��P�4�u��n��K��7Z�pf	�����oda�ˢ^��l��I�3��~p�D��יÏs�QB��2��x�>�):mA9���޶����v�7N�i��ܭ�4M���#��j��T��*e}*�g-�('9ֶ1��7�0�;h6aW����H���u8�y��P���Iv[�`�<r(-7?>|}��ڜ� �����$�ײ��^�S1H���x�%��x"��O��G=�����xˊ��R����e�8�8���=)L�QF�k�x�[q�"hyP�o��"��ͯL]�H�SRt�m$�ѧ���GGd��f�Bl$�B+��o(��3�pgp|E�"*s���/�ػ�F��⛧��@x��:]��u|�p;��9�p�a�e�Y���Z�z��3��|��{)�r~(���3������g֎���_�m"��o\�W��2>!\z�H ��#�-3�F�x+�/�� �"�}H4�_-Ж�p���Y1����&֙d�s OS��H#�;g�d��kB"�]���tO҃�J]�/��_㒡~��E9���G�5I�(
u4��������~�����K'�����f�)g`�N��W&�$lV9�>t�' ����轆��\�91�R��[Ҧ{&�͗��݂�V�A�m����*�v����%w���p�#WW�+�VDk~k��u��F�<q�w�c����������7�n�?Gj��qny۰HaB�f{k-VaFw�\z2P�Ed)V`�s̎�8�>� �\�gj`�A��Y�&�"ӷ����iVG��if�ϱ�h�(��^K)G4ާn�҂��1��Eد	�Q�'�\v����Te�Ո��pn�y
��.�e��G_8E�I$�Z��&5��a�&