XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t#��)��!pf.��S���0�B][�ە#�T���a7/?yh���F�y@8����S	4áК�(ӆf�ƺg�X�Xk؉˙%mr�k�f'/y��R�*p��j�f|���F���~λ����Cý5-b�m���������GA*�k�)v<:Df0h9mAT�>l����/��s�r5b��-o�k���)�w��k5c��gOSSq^'|:Q�����=uh:/~N$7M���̒�m���tNU����{c�Q���iZ�D�Z:�f��w޻���^�#��j�^����\��pZ��X���C;	����?R1�#��l2M,?rBJ$R��`y^��SԄ�o&��}q_Em���q�K�������X;�*�.���#�Q��{R���g��B�6��Y��]K�b����H��_&1s6aaB����e�'�^K�\�IF�S�V�r��[�X#SD��1 �DPۤ�<���1~A?MZ���F��L3���P���rT{P�l|)��C�eX��"� �x��:�8��yc�%hJ��Ҝ�"عmQ�Kۋ�)>��"�7���H<Yb����9!��
�n��u�:�-�a��zZ���t/��\+��A�w�S��-�4,��q$9k�lI�+�2�2f  Z*/�R��1[����"��J��������rǴoF��L������JG'����;�d*5l�jņ�*��]w����]�����-����D��B���4���^�;��<XlxVHYEB    152e     580{�4�ޜB��it�\G=B*�����O���i ����/��!�T�e��H�Z`�ض��f��&b��Y��:�,RN������T��e�)g������ �����YYo�l�{�%Pʪ�ٰ��t~q{cr>&8����	�	�.��ԷA-�/��?ph�v�{�R��e�E��Y!���*̦J��9G��$�� ����(o����W��[��'�W��q�2��M1s��h%���[]f�:'����=���1��!+/4µݯ�ϲ4v�Z9��77w�����.�Y���8�mP��l�f	�\[�A*RX�P�7W8�~����~��Z�8�&OW��/�F���U룟�
o��l.r03�\�y�S���B"g��W�U���R�I!6����(�y6���-$S��旼=���&n����1����3ܗ�ߩi��0.tcѺ\�°����R�x�Y�c��嗫�	}! �m���\�[{כűԶQ!�lB�:b�cpKܜ���a�*�� ?eY��.ߚV��//9�E��u�w��ϋ�0�w	��^��A[�HlS�&����(����̍w�.bE����s_�ʦ�a�RƥЫ�̢�2��o�e�y+�� P�wz)�T��u�����@gD�'�l���Ai���Qb� o*�e��86�"�s�X7�wgZw�� ���V���������{=���ŝ�ʡ1xh`ݵ5i狥�@<3�`2�m�5ʽ?���=帡8G~l���@�O]��47�����\�DV"x6�
��-�f8V�(���ڬά@�xWr�s6��-rz��]БQ�0��m!�x�!�쿪@P����/sU��k�U(�t��!�l"�ü\|�Q�D�����G����+��\�ǂ��t���3��f�u�?RP�HT(�V͞c�ذ����0��q1p`�����%�ml{�����iTd]�(q�,�د
�~pe�,6(TggIE�^b+�xŏ� �lp0�=��F9��� s�J�~a$�QƁ�}��ԗݎ  ��9ףp�Zģi�=A>�^�:4���o�gI�xQp\���7"��ay�i��J�V2�g~,>��䯂ū�*N��\��1��� �z�	d����r�~q�X���� �����72]q����q��`@1ТS�r�w�P�=�!��5�Iӧ���{�Oo��(��f���v��8ﮤ,�JU@7�Ѭu��i�S_Y4I(�ླQ���bi-	�尖qN�P����'�1��`�����tW��!����"�7��%V]n�q�w2�k�f6,��y}t�y8��B烓���z�D��?�&�}Z$I`&�&�1)���Iy��()^�h���ĭ$Uǆ��rb��3��N��b��J�<_�PJx