XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^�m���*b	�����(�~@�>��!�0�=Y1C�b��]уJ�}ސ��t�. � ��H��	|!��sE�y]EN���?ڥ����ZH���~�T� |W���:n{�+����ٟ<���d�s��Og0�I<���*����Eie��f��Ǝ= ��=yZ|�ދ�x�	q@|��{/~��Kf���s��:�
���!��+<Esf��Ց��ȼ5y^�bj��e���'l��Y��;5��ٰ����5������EEk<���Z��}y(�Ԇ����� �t����b�+m���7 �s�h�X�~%>�(�a`���)�.J��+���mC�*�MOY�f҄!FK&"�s�޲��'�*�b�T�m�ַ�<P��jh4�D��0�L�侤�>!fq[�y
1�64�1�y.{������h�VD�`��k�܏3{%#���NVy";e�2��լ�_���yj]&��|g�32P��0�?}>c+9�􂠂��xY��t�r�|Bm���cF����#�3)�rp���)� $�C�6AƮy�e_%������3�,	�X쫿R-.DxTK�0�F�X��iZ'�۞���=�"��Y�f�#�H=�����
 �Ky:}hٺf�_��d�S���B�P�
�h�N�h����Y�h$O�%4�!6���B&:��@WS���'�5��U]�[?�5�!$IE�H}�^ӴZ�k=[����S�cM@V�~gb���7O׈ҭ�XlxVHYEB     ab5     420t�HfWq�w�9%dm很l� r p2Xv�������W�$:��_�IxFY����\���f"�R�/Ÿ���f��πO̶������\}��6�N�?`�qL�|��H�|hh�0�,�e������	o���,K2�}?�}F[�)�f)���7q��(������|���n�Օ�ѵ��*7F��s �i��v��3q>��؟�1���������,�'�zbr��})���T�! ���c~����d� ����k�F��j���>���߃l��i(���XLsվMS`�q���$�I��址�,�l��u��K����e����'�8�r9L'�/��H}<S� ƷM����lT��KS�~�6H��j�\%v8K"$���GO]����J���&W�ыCd�����]�3����L����"=g�<$�>�.���϶�1H���e*��[W�B���y����	���	�<0�ƭ�YJ���`�Tv�8h��#��b(׷�Zr����A#7�W�� �9=��a����~�
|��8T���!���F�[�S�8�(	��;G؍$ZO���	V����z�n�T9+��iOy��"�Y�u�-�;�bD��*_��"N/J�A������rdz����:X���u ^��&h�3ÜpX�
�!�����JV��=�&�v'��7Ұp�z�h#+���G��uE�|�̡3�{�;ӵ�	N�r�d�mo���~0�~��ܤ,�u��BF��b-�1��9�Y����ġ7�0<a�;�%��l�Ru�(L�6�^;�a���X�#+U�:@Q�� f+yo.5�ڐ�r���Y�xQܻ�w�6�*��ޕ�ҏ�u�\A8��c��� f�4�^��*���K�������S��]1�|CP����/R�T�5�UM����x��#=�������[4>�����:����]�	m�m|ԙ �ITO�m���kOz%rHq�K-`ǖp����Q���� v|�z�e$�}��9꣗!�*�ro�FnO"�Fc�&�L&��g-1�