XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#m%��J��_O?��A�����#��!UƔv�@N�2y����V��	=2#�n�#�R����t���,�P�����Lx�L�3�7����b�A��-��Ї��HOGw���w��e)��U��DWj�̊�x�6Z�i�sl�����Ǳ%,`�鏤\"UV+FtQp�B�=�⇾���(�W��dܤn��X�/��L8�Ч��z�/�g�a��`�,���V~�i��9#��V?iW�D�-��Cc�ʩ�7�y{��o Mp�XG�	S*�L��6S`��w\h�K���S�!1�"a�G=�£��!���׭�z���Q��q��m<��r"�
�7�U����>��F�����<��W�����	!���-n�d������2"5����k�K�d���$�����P�������������Ď�����E�T���`:�r?�Xr������/
�hˁG;�B�>������4r�n��/�)�"����fx'�ƫ'���g���]ˡɭx����.-	�7��Ԙv�I�uD*��s���}�PE,�V�D�Z,��ܠ����z��A���*�� 8��/����x>:L�#��󷿥	%,Tp��3�.�K��
���x����8u��K�u-ta�l) ��x�l�3��H�끅ܷM��&�B�&].	Jt�"�;ֆ��%�p��\:&O�[�W��3|��{��N�.X�+[�����7eh������<XlxVHYEB    2864     8d0��y�$hu�̢	���Mn�S�:����_[��NH�76	�]@�2,c����R�������8���?�C��(3�x.���>��A̛������z��o�KZX�5&��냁��u	���Y��#<��cz���!֎oW�pJ�@r9��M-X�bZIy�В�Ni�Fm����2�P�֠��6��X�P�)��n���ٞe?UQ�#%��G6]�\|�N���,��ATO����F*l�jGʂ�kF+�j��x[�=_��G����u�NŃ�fl�S����{k��f�/|<#/�~���Ԏ�Q�!k���|����	Hp�^��� H���X!4܊�Zԛ6~��3!q�
��ܖq(~�I#�ھ�%P��S�X=w�g�tz��t�z����T�G&��MU�Z�G��2���x��k�o�;v�G<}��b�z�\C�t	f �)�p��8��·�Sm�h�����\��?�Èz�����hk���J�� L����x���ֶ؞��i5W��m��"ACa<�����ygL�x����	=������Y���;��5$�l�X(=�Ԩ�ya��a�,/oҽ�ס8t���U�I\1F�����B4"�;��6M&nKҩ� �K&(�(ק��G.��K�zj�%7�di��*���&�����0�����E�lY�O� 6Ln֪�(���\����A(8W;>+���N٬;qߙ"S��T��a�MeP���C��)�s��|�5��r�^8��V{W���E<�k嘌i�7F���n<�`Q���:�A�����ty���O��{���D9����E�qa�ù��Ɏ[����%�8�=��"���fA�J���U��o�T?��{��j��=f�seT{���&V��͆\�Rc��D*n�>�"O��Ӽ�`<�w�U�j�Z,�l����/e|9;���92�7,��X&�	�)x���C^���G&�!���p�3u��a�s�lA~�N���`�j�E2�"�Q�
�������r�2�FU���O,��e�%�qinJ"pU����w��<�m�_�|��'N@�6A��փ�W����#>@@�<Fa�[O3� ���5u�Q�-f]*�,R�l���Mj��うQ%�Z �4�Z���E��b�n�S}�5�������5� ݺ�)n𑅎嶐3zӴtZ��*�(��Y�_Y���)�p8T B�w���u�;8���Nk]�l���wE�M�_ܲ��T<�aN�m��f�2�}�� �pp&���	�O}>_��%y�4�O6�Q/�Pͮ�WdhE$�SP����jb��(�\���&I�Ϛm,ߏ��8�$��E�@,�4 x��L��@|==+�S@�]s��A�C෭����S��|�	8-��N�!�6U/vN�Okcs�x��+4�����d~M&��>�L������g�{�讂g!ܘ:ﱊ�'����Y������� ��kN�e6����y͹�ǲ�T�!s��4�$�P��S��Z�t(���.K3�mmP�/k珠#BDt�<���Y�2#hb���y���4 �ؚ޴�˜;�����TM)��
i�`t�����������)9 t�k�V� _m���������=�n4�T*����yl&��W�>H�+C�������H��{
��v�v�҂�c��j���f7ñd
��i�S�V>�v�۾�(��=)]�@�U��s>�,ƥ�il�V��N�R�U9�|3�"��0+���A'��;�:x��
�������e@�_��Tp4�K�d��գ3��v)ק��-pn�e�hA�Rԛ��T�x]A�����I#g�9a���.>,��>�N���#�0�N�	�������b.����H�w�i�z�h��N�b�2�� �nCy���Ui3�5Y�<����]/ɽz���o&�Y�#~�.fꔥp0�(�{>���F�{�X>tvz�Eo�0uY��s龫���8�]��]CGC�*��Tf�	�lt�Ma�#�9���ļ3�av�	!X ?M�qw
�����=�;� Hٻwm�,�����s/ͽ���QΓ�mU�?�W'�U�,���&CT!�֕-d5�{@Y
}ڸ����R�4��9�ۺ��g>���z�������r�zȘ������AE9*�2�sم�P������~�>�XǺ��T��H�T�﷼�7���