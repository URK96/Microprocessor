XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%W�Fl�`�\:�Z���ذ�,�Һ���e���ct���6<H��]����]�,$y��j�b���[[ʒQɜ��� q���bӊ�����>��BlS��\���H�å �s�z�P�#d�b�C~w�h�hg�2���i�ۃ��t���o;���C�Gѫz+��u���P�O"�P��R�&I����̚��f���E���Uar�nd�m�����	;�-C�Q ��Ƥ���u@�F̾����8q�Y�+б�Ei�/��rw�U�< �ť82k�nU�k�q������?|S��`�e7�͡G-�w�έ�5�n)%����P�^bu.n�x��K��h7�;�7z���Z�ԥ��,a$�Z��ק��u����TK�>x���}j�}q����1'Pl��p��ϽN���173�E�&Y�m���/�[�L� �w��a�0݉"��������T�>XKe�:�*�h�G6�G�A���=��v[�pb��"d���fj0��nXв���#�!��m��l4)�_2Z�c�CE�&\�1A�^OL:9&".t0�2�䚖3ie�Z/��n-GF�̶���351��U�\�|9%'�9�p�@���'�9���6�+E-��Cs� ���ǇdC�t<��*̘���Vne[���y��-�c�19��΢�X�d�;ύe��� GQ�j�h���VO��n'Zא�k�k=��[�k*���&���i�{�zն=�����C�Ct���K�k�XlxVHYEB    1d52     7b0ǔ�����Q�
��њ���DZṩX��dv�HR�h���O�HDU��$���x#�H�ߺ�7�ڑ8����ܸ��k���J��I�[�y������ş��βHG�h�I��4��w��������J�FW�R����ԍ��>S�n,
cߖ{ܯ	d���:"\aHoM��&_R�� m���}'�֊�HN��/�+'�D��ƐJx	��h ������s0�7���C�����P��^�e���@�_�6u���u��z��X�J�xmE�N.n�[;M���}~ ~^}�$i��DIis.�t	���9Y�U�X^Ԫ���SG͆�J�e&[;����5v��eK9�0G@z�����dlD�(K�%�A��)���S�/���S����ι5%�FN*b�_�2�@ �pt���н������PS0��A�$`_Ϥ��9����������M}I�|���_3��B`sk��	;T��Ě�b�%9�O��k�R��
(����飄��\��} lO���Aqބĉ��v �y����̜8�O�����]̴�8����Ȉ�l�����w���5;uw����IU�p;Հ�D6N��G?DQ
y����SVs&�` <�l�D�����G"����6ω� Qб=�آ,�u����4�d$���_��@5GSfI{c�&`���G�iZ;��L�zL ��MX���NZ��5��G`S����vL��J����z��������ݓ�vh�6_��. )���1���?P�D�����N�j(��>�T�t$���z��-�3��
�7,q5L���1z����>Qfcb��v芷� �IpZC)�>��KwS��m�WS�X�dץ��#D`٤��H�!�� :�i�
�`���Q���.�oͩ�XX�|��n�`u�󎊆�$�mY\+��A�,��j���c<ؕH:b�@��e��X���Rc)�i;���й��!*Y�����uk����h�ܺ\Ix��|Ԧ2��,%
�Lw��S�s�'�+�^���j'���|���<�H{�@-�U�j���,+����J���mJC؜91���<C�������� ,ѧ�S�SVv�ͻ�?<���z�|�|�f;f!88G����C���WG�;J ��JkU���7�Լ�,�a=�z��GEJ}��$�GG���T��;O/oˮ(����'ݛ���X�h������:����ś4	h�B<�+��i�a�d�\�*��
4b�)�@f%����!��d$=�U�V�9�<`7Zǚ	���W(�y��:�x�t�{gN��~�o��!��mD�^s~�e�t'S�%|�LF񡊣s۰�)��Մt�?�.Z�l��S��d}$�;�ß�5_׆ҹ��
�MU��?$�=?3��(�C���[~�t��+yiJ	�R��s�q�T� �I&-P5�.�e4�q����p�2��Qzk?�aP����Js�/��	�7Ll{4h��=-]��=��&<�Gia��pcP;�&�$
K���7GY����oYװ�S3���v�֙9Ǒ�0��w���Q�V�"�t� �4�Ql�Vj���df�܌��b���ST�Ѐ���bHZ��ޣ�1���7g����0�6Z�d	�(9�� 5�	\V���`7IDl|]�J!���mmw�½��/�`�2C�&�Ԥ��<��<x��E�ޥ+?d�?�w�)Y���6�g����wgt�2��4I	���1��O��ɓz����e���:����3Θ3�%��6%Q�,���'N�7^��lA�������u�NsX��ugׅ������z��u��\�J@�����z2�2{�]�����6'փ�Êz�y��
[���k���1eB(��b��5��MH9��m;a�W�/�2� ��y��������G�������Tڷ"��t�I