XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q���Rj�g��+����5�x޲o��9���h�L1��5>��'~"�1}P������3����J*nF7��-$�������"��Ϫ��i���c����;��=\ry�x����Yt��L���j'#��g��!�$H�������J�C8B��VM�Þ�S��F��ׯ�S�O8�?�;�W��������,;=X ��{�IU �:�I>��9W�N��?3F��G5�f$���^���rd���?%�FiuHi�#�w����}w5���5St܉�3E���,�xK�TE-�Xh����e#� 
��%o��)�;~E�_](�s�ՊK�Q+�UG���?�J��vW\MfX@;wUȴ�h��*�-����'�ߩ3��Y<(v����(	d![�Җ�n������-*%u-���ŧ�y�6K�M*�G� _4��{��_�.�V���{#��x <86�p�T��f����q:#M�� -�b�
ۧ��[��y��`���?��&\
6�����L�9Cq�)`�����D�J�M�ڣ���	�ɂ"pp���,#�6[�7pY��/aW�O���ny]����I�0��VLh�&�ލ�V�� �N2Y>�S��3���?1�2��
|.�YF�h�s�s%���C7���|�L���K���l�G��J{�U�EE�U|�ψ��Fƭ�^Ǹ�Ksi���6Q��MK�������D湉�jO����vm��x�����~�8�Y��w�A�m���s���ʕ�XlxVHYEB    4d93     cb0�ַp ���c`�֋QO�NE"�+4]�O�˳���P��,������	+���\�B)8hFHH�Jg&3��~VC.�`5W�L�c�L�\I�r� ֋K����ö�����+/˟˛�6��Zid}���<�D���ș �>�D�D{�����yȚ�zРAˢ�P�T��=-�D�,%�;؟$�7D0��raA���f ���u|��z.��T���� ���\���;$���$jq�h<�=GgΫ�����魦�L��m��q	��Ȗi+�sv��Oz_�L��c�����J[�1�ݎqC|�N��bҽ������S�r�A!W�K����E��X����}-�p�q��UM�aa�bV��sW�pq"n�Ė\S"2۲7q��C�Fd�I����@&g�
�T5F�5¿��7Oononׂʸ(�mr�G���Rp��+cN*�Ao	{�dfךf���f�Gu�����va/:���V�U,QY<H����&��^f��V��9�1�D���zh��{���M�	I�[U~o��g�c�ԛ"d�#�w=S>�y�Te��컸T~Z��==�j�a��:�x�����z�3,�����~�g��i��we펄�ߧM��W�z����!��ӑ�؈=h�>�[�	U
V��OZ���%ϚU2y^X:V������q���J-`+$�g���Lġs�{}��m�e~8�y�T�_��!'D��˄��P����6��L��#7)-�;�FPv�����v��iXǁꖯQO��<�0�ry���}��ܻ0l �	
�<�:b6�æ�]k�x��r��_�4	IN�n���s�o(�iL����mh�Ё�fL&�����n5L��HzM�����I����j�<�	�5���:�X3�+{����%5n%;���zyL;n�^o���`�x���m ���/	���d*i�Ӽ�2�"p�!�K=|8F;N�}pn��O��c��z}�tdX�������r~����,��3[ҥLB��u�e:wο� ��+�y>��*�K�/<'�au�LG�D�㏪�AQN�S>w�Q��W4~ {�6��m���v����tQ�3��n��KH��!�}ڗ�
3���|�z�(��Z0\�?J��s
�s����Y,8��}��g�>�o���h�P뗨��ߙWTS�Ѹ��%���6���6�z|7�Kϟ#K�[`����)�!^�"i3jI�M���2n�A�K�	�5c�G����s)E�c|,_�I?'6���8R��r��e��)���+5T��MTM��Y�Zq���z���;w�)�ҙ@R��.�'@��5�d�7Zw����V�����SZ �	H�Ő���X��@�EFP����'����(�8܌�O��Z1�5������#�._|!�z+��2F�翏-�U�8��p�q�~���q2^x����j��Ԑ�HԌ�'�d�㜘k��dS�/���g����/y��ڡ�4���A�(J�Y$�(��%D2��R����d��˅w�6�{Az0�����d]!:��T���I���|���0c& ��=Zss9�]4�(W;��Řa�e�h���@�N���'
�f%��mP����s��w�|�u����܎�Q��'5�f��R���	�e'�����2�~��bR�*U�H=Wk5݁6��"@�h�+<"@^s>�蝞
&+���!`3gI���aBā:$���uU	�
�N�6�/��V0�j[#!�0\�ʕA�cv�;�o�	߿��uw��ǋ8�4?jkK�g�<��r��]����Rf j��o���o�� ���x��*%�[Z��F찥��x�*e	�m�p�"�% ����Q�|����/��'�`���N\+�k
���������Q���|��Q��U�7�� �P��!k��(��c����n��b�#H�e,����xJ7g��Oё6 )@&:��ډ����7�{X��[��m\��8�!�@x����)�*G�:oQ��~�b����E��U��ʪ�K���m[��Y{�vM�l�܇��`��4�+�,)V�T�K�}���<�����lƁ@��w"F�'36=EX���rH�A���>p,��H�,� ���>s[ܪh %b;aധo�}�J�Zs߀I�-%lhя*56��5 ���_rq�DP�욷 7��b��p� �I�pTS#՝�+%���.��Z��O�7�O��DY�s�<N��xK����&��T�p���_�����M��bg4�.�(!��C)i;��jHi�Q*��Y���@;���h�(���tEf�]ȀIeĸ��Y��^�����EH,�]S��- }[�W;ua���)v�>b��'l��|`r��U�k9�#�E������ZI�P�c�.�lؼ��*�n:�T�����kag��x��J|�Q�2&��+�qF�W��t�3d�̜&#Y�X��33}z!]�mj�4i��j�&�9KUi�l�{b]F&w������S~b��΅/yB��$�_��%�R�؉�����׳峆)H�{|b��l�֕���R�������JeH�\�W��I�I�5KХ���y:	�楇����gU�lX�akDl�D�6J{� V��a��x��`���^�`w ��PP�-C!s	+��e0�t���Α���C#�w�X5fe�XX����J�a�V� X���ӥe^g���;~�SDű���+������pP�P�(��{0�d�?��*�5>���9��������Gӵ)�4�C�\Y���X����s`|I�N�̛�|ۚ�UL"�.�|�p��R�YM>Kh�w?J�J|u%�[��B�Ԥ�b�DR�AF����S���<Q1�^M�p ឋ�0Ѥ|85�i�I���$����Pf��N��e�ҏ!��ؑl�}�A����_���꧛�uK�U.� JlV�F]�X�i^���Q�RO��l���L"*�L��� ���Q{nN�Tޢ�Ң��G���c=\2��ܷ�B��av7�c&�\��9��`�F��O�G^}��KG"k=� ��}{n�/�fl/Єu�ܱ�j�j�FTE��B�H�RH��.��P)�1��ٞ/���+���|�¸�r3| �B�$�j�B�>�}���ay-��Fɫ�C�Su