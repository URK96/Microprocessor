XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���q@&w	st{��/�0}�ml�j���uN�2�Sf��u�P��(��x��󕕋wP)�ݍN�͈'IMW��@ޑ��*��G����E+�c0�C�K����K]˦�h���qU/���CG�/Q�+"3��cX�M�~��P��@	ڧ��� �#��Y�gVîc<�i�����禫����|~��Dy��
��^o���1��B'�#L�X.�E��ig�$c�q�V�4���_�Y�k:nM�C���U�b)<4�<�ݰ��,�Ii"���Vc��.�%n��E%<F�(�g�{n:յ����ș<Q�u�+z��G��֪��>�OA�Y�����-�V�f�~F:� ?Pq����َܽ�uU�Ӝ/,�tݎ��i�����΀+TRAd�]W��K`��o?7\�"<1y���l�GX�\��q��tC>h��EՇ(y���=��� ����:��Q����q�o7H���p��;$�,�J���c����I+�.�D��N6��@n^?��1��L�e�K�i���<cཚB��Q�A;}8�>��KP%13܈Y��UV����C̏����������YQ���r�/i7綝�C%K�6��^e�.0jp"N��5ᥦ�T2(U1�9� u�B��
���TՒ�N[��hB��y+��Puy@rfƥ�_�aa�.8�W��d�Q���_������*���]5���.>�۳�`W�]�����!,�h��H����r��Wiv��_��ݲ ܃XlxVHYEB    1569     590�qx +���E�(e�ͮ�)/��K�Cߊj��L�j�z���0u;i3K�>&���4�Э:�<=�h��n2�
s���Y>�=tS(	�7���f�'�  ��c�1#z/p��J�G�_�@�_�ϏQ��"o?4Z�¼�5Z��{�h�W�h��N���l������}e�e��ɟ�6���鷫 jt����q`�ۥZ7ź�1i�G�擆�%G��8��(��E��h]D�4�4x
�q6��F����T�3P�S�����~��aY3ц�J�	/��t�nE�c��i���@���"���1�r�:4��p�I��T�U��)��\��h������g �w�0��k�3��d.4Z�2�8�I��8٬��|���l$�)��ѕ��5�·);�  Q�#��)�������p!��\{ e�N�A���D�V�E��n��o?��23h��/�7�I�
�{#�'�§~
����u6x͒	��Q1�YG�kB� èrfg)��������uY&ʌ��\���`;��#�����7�++����M��D�ѣ�#�1�pn��xrԖ��f<�	(�9_4�(V��?R���QԌ|��⹸t�8��)x̹8�+�~X�!6����ѯLbM�9�@��\�Vs��! V�$ G��-��_�!�t��� ��M�qA���ff�95�
bs�R��j���IX��"��O*����F�.�3|G�0:ٍ��_���YKg�ƫ���8�gupn�,	e��E��z}ꥣ?�>{=Ř�|�
#�x��!�6s ��(f���D�`�<Mx�eYdʛ����/5����F����J��1��eR
@Q��Z�W6g ����+ȕ�u0�V����D���%��[($՚k2W{�����j�o��9��T�/�ɖ{C�fε�`x�����=�]1 �%���{WXR����^��\���b�)�'�ñ��*�K!Y3@^gk��F�=��b|�U�}=}�kxp��LV)m�5�G�W|�?C�lI+���E�b�^:s��v^�6,ˁݭ�OW���7��i*t���ͩ�נ&����1߉T��+�y a4]_�3�3ud7V)4d���ϣ�qe�fD�;ۻ����&�t�?=]���/�:D�.7�i��+�@ϋSnvv��#��k�'b$��� ��,Ў�
��+��� �&�Ix�J�0��'i7Z�J�� ���1|;t{�CQ�`�%�[?���j5o*! n�Ql�{+�U@y�i!�A�:5(��V�P��!�%X���E�W�L����x�����[X�N¼aȐ�nF��1����=��H�&M�Fx`��������2'�6�!���s	��Z�-���\�"�������'B�F������,�ڮm��`��|��=�:s�B�ȅQR