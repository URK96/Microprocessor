XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.���ۼ˹؞�_9�;��\�W�>���LgA�7�SUjG��zRɫ%�.���Ә�Q8�HZ�W��uY�$���8�؋>�����|��$)����SO(�`]� )G�^�f�~���]�����ܷ �l�Ǧ�7�2T��O���]ud�Z�)�R䙅ʗY��x���7���<���1�x4��Qˮ=��LM2��Ɉ�(���t�w��C�oa�ݓ�^<�3��[�p�R�q�ɿ�d�����B�`�x����{3�&'Ϸ�7��Q�ֵЂF��ŋ�uI�e�O*qa������>��Q��������G��~r��l'��7��m4΄����g�f�@�����Qڦ[o/�8�{�X���B�tK��*34�~��Z���%��'{Skݨs�@  
vK�$VсD��L{�d�I����_��A�{1L/���<+���X����9��6�����6�ev�,F6!��'���JG8!'���X�c��u��0^���ux��d�H/�s�!G��m��C�A�at!�fCs=$وs�r��|���C��*�F8��KQq�+9�[�n��c�78���.>�w�:~~�Y�B�#?mA�!�n�]o�i��w�����Z�`�Q�S
�p�J�
��+���L�Ҏ�:��O��4p�5̐�
H%���"16M�K����W�]���A��ӝFV�m������;	�J�@��ڥ9f)0��8�ʘ]0�S[$8�u)�jC�R!R��?�|3a>����qN��XlxVHYEB    156b     590�egr��^���L��t{ޭ�W:	8e)M�̺���S��#�s)�T'_�2|�R��P���h;�`��C����B��+�#��&o %_&
r��(��(�Y�.E��_��
}'UQ���)�{A���+���*�*j�-Rs���e,!�k��P<��x̀��K`�"��=hzf��#�ȺR�����Υ���W���
o�Y�����D[f�_��`�dGx�͡Q������'��a���jT�$g�L|�(�!�/6���&P�Duf]?A�X3 K���e�a�*0�{�u��O���9�3����w���h�j.ڄl'�n�e� �#I�r}^gϪY�B/������d�,��L��g��#^��Ý�,��f����8��Ï��e�9Z��2���`�>M��7r�ܾ��^f�m`�Z�����!|��uB_k$�\m%b� 5�9m��m9�^V(cI}�L��ӢV8������ƕ�^�Y"���{�SV�Z���w����э��	wn��|#�j�T'�f��B)q�0�*���ZzW�t=�"�Q�"o�~���u�ϵ�E@Gw�<���~<!%Q8z�b��76��"�������^���	�\�Z:��eo"g�]��f�ջ�ʹ�z�>�(�{@�bw��q�Gm�5�����Nf�B���@� �k�wk6�g��i9��9~ȺT��.�ԙ��z�v�.���R�v���ꃘHKZ��01��P�՘|1��z��UoҢO8��`򵛣fW��aa�\��."౿힇*P1��T����hO�8[>F��94a������P�[�fVqr�A�hE(䜈kJ;LLKhV�EXƤ�T1�h���ԏ�w�~jqa�}W���F`�9^F��-6��.�c�`ŋֵ�.Tա���U�!6&9��~�!3~b?Kh�íկ���g�g�\OaAN��p㛭t��ӶE���ە�X}Oތ�;�"�cDL:C(~�@b۰V��;@[_Ƅ �E��XK_c ;�W���RЀ���.H
��6�̖V!��G����c����$����kw}J�����BF��m*k���ϴ��	���Μ��TM��u$S��G��i|��M\��I���t�N�+��\tQY��v���RT���o�2����ȅ�wî�3�\؎�5/�ʿ�(j��s����gJ�|�9�
����N<�s93�MKwT���
�����d|�̙[�H��V���)O#��U�e�?�olH�b�{���\cͽ����a3�w�_mz��+u�0����4DB9%��n�/���:U���M�4L��w��i�/m��p-��j��q�*�.\�\6�cL��/e��vo�˙&�ֳ� �����6'ĉ.��@~U�t�����L,�ڿ�0~�&��