XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��N/z9'|����c��V&D���[�s�1��9�Cu��D�^�h� W��p��5��@��^���Y`-#Lq�e����%����Ѥ�i�|`8��B	s��ԇ^�c^��t�
��_���j�u�/�:\�C�� [b����)ޔۊH�o%ͼ�x,6��}�,P�=�������������}Q��I���z`v~a�au�Ҷ�*�?��c�$;$$g]�|{�`������}{LFA���	�U�pթ�sOaٓ��oB�ytzf��!ƶn�X�͠0�m�oh��j�zr�JD!��HN����%�t+<j�@�A�E��z|r��# S�?�"�_@��|�;	a�*��I�����"Ձ^��Xo<�� ���/�[��ż�z�E�M�N˭�Ri^���N ����G���j_�1'�v&��z�ݥ�C�V�n�Q�q�Y�n�C@�چ�6'vģF�¸k�?��R��O�q�V���H�D����Y.�Ak��\]�HH�k�+K�r�c�#h����̻S�v%���c�2��/�*F��-k���4X��}ﾔ�sς��h�����W�εS�����9G[�!��#�� �zT�ϵ6*�2P��6<���xH@�δ�Q��:��,�T51Ŭ�cJ���]+y-���Trj����q�l�RC�����ƶ�"42�͜W,RO��Gs�F���\}A��kt���Ѧ�]R�Ą��6�xk�rƯ�\D�O���=v|�{�@Aj�R������3����>���m��J�4XlxVHYEB    1cf8     790�v��zT^���)W����-U�m��z�Ox��>�y��� ��!�<���yo�]ƺɄ���A����ǏWu4(FFޓȮ��?�|+5��gU�)�V�, V����uOI�T:^7�8j��r��/f�;��90;l��K��VL���T��(���~C"H~�̜�f͎J}TWձ\l����٥��A�����# v��t���1��<M��Y��f"�E��u��
��~��+Уo`b�����"g�6����#�X~�z��@�`uK(��H9�v�rjTw����{��A���P��c�0��II=�l(1o3��=��r��B��R�]/��T\PU2<�|����C�${(C���r�=��?:�HeZ���p<�.&�>`��iHn:�]����5$��翅a�a�>�ͿM��)���#wU��O��v.�ޔ�I��'	�_5!>t�\���S�X�%��)� G-wM��I2!����+l�+u��t�3�pR���;����uk�cP����T�s���`3 ~���{W�\�j�#�0�f'�"["�y���ڽ�d��l�=х(&@�|Ibہ� �$�
代g�T��>�F����wj�}(Yȃ����-[.C��#�.f���0�<���<��T}+L��l�����=��}s�r��se��N�_ �Qf�S��c���*���_D�;W��@'֘��]j��:�j��ϊ:�;�����0��?3�J�8�o���NC뮄�:��mկ(:)H�
�L�J�Ӟ�)�$�W���ب����K$@
Q�JF��A�z��"���i��[�<+WA�_�Q�d~�����a�2��,XI�����~�vh8�Bl��Y��C�˔A�=�\����P�A�\f>;ߵ�{�BȁQ|� �S"��̢�"�1�ZϢK�8*�=^��Eqj 8�� �2�K��@b����'���& �S�/�^���;SX��(DC���2��*�g���<�CSe9_�l}��݄�DT��1�W?u�A�tcE'o|�-��e/�Jqsㄡ��[v�G��V� C�d�q��5ߺo�G��w�8��T�b�"���g���/!!)��.�p]O"��_�ʅ�>�M}-����O���ۖ��5�/2��/���P�x��|���w��=9�$���)P�ϻ�����N�^�9��v�dY`���D�E�~Eݑ?���50�����Ե�	dl����c��$�Y0y�tư;��J�_%�$�AY�.��m=lu�+��7��v��[!�gUJ&���:S�J�pǊֱ��,��NIB�¤Bq�>�۴L��;�9[y��bu]�9�ؒ���l��(̙l��yW"0,���8c�0o%��Lӝ��'̖w0"Q�˅R�R�n��y�B~���)�8.���Ւ��f����2�33<�g�&�� �d�����?C,(�E��1� ��h\]��;�<~l$��7��,ډRp-�͓J7B�Ӄ,BR4y&j#�E��
��]�F�M�@�yYY'��.�i��y��c�����`����Q��<���\\�	�e��R=Go<RV�Go�]�Z���x<�g����G��0��@����s���%q&�u�e�^3 �BǮ<�5yԌp�V�.݋n�N��Te��yPb8�!U��Z���B.��~^z���W��|���w �����JR����o���ڐ(2+��ɮ��x� ����~�X����PA�TJ�Ja�թ��o�1�$G��x�O4ke�	71u���.��W�+��6���� et$�bg�6���n#�rb����D�!�L���<{�ۈ�U��Q��n�P���-RާǶK�"D����ߢ:��4�w9\23YM��z_�`��T�t�����r��