XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��َ��!�׽�R4%Y߳����2td�`V*ucj~8����;O���G{��:����=79,ۤ+,d��wMި�[���j��o�b�6��L�;}J�%+��wB��	�u{�a���.���Z}&������6)�ehד�*jy�x��%�y�<�b��/6��"���RH�%:�7�ƫ��BR�2a�3����<�;�OY�/\n�e������ZW��
`��bH�� ;�̌Ǌn�������IuF�~���t~��(������h	&.艠]/d�Ցz
J`ha����ǻT�j����On9�~�4	D�]q=����B�ۘ�����o?~=CuҬ,OU�v5��Z�g��?���^��Hc��~�SF6==˹���͖�Z���]��.P,���1�ʉS���Zy�P�Q��a44r)s���B����
���*���F�,��Lu��}_�{~7��(�]5� 7�r��o� �;�-S�b|��<ң�{��_�_�McPW�[M�]<|��)�i�M0��1\uq�"
�<R�V?��o�ԸI��$�yB���O�a��n�oڣ\�U}%��+Fr�[;�b�z�N��?A{U`R����[{k唨�P�{~0aw_�[*�b��O�r*/؀�l<��J�:�\U�d�Ǽ@�Д��[T9ޜ͂4�d����l�j�w�8>�S��qq�±��A���Q�t�O��\�ȫ?��?�ї�T���[Ђ���[���'�:kȉǉ���Q�yXlxVHYEB    5ff3    1040£.�[C��N뀩>�-�_�o/���1[�-�kym�,A侫�ݭ���5�T'k*�5W��`T�Md��<�:�m5!����R#E���y	���o���h��~�Ȟ7>�ޮ{�j!Ҭ;��6yk�H;���l�x>��XO��>|�����9d�����2$��M=5spu��c��\}ʁ�5S���F�	PI��m�;��bũV���B.}p��}8���ģ̾TN t9r�o��x�|W&ֆ�3��65P���[r�d� w�BG'e�E���૪�@ښ�b�M�.ݛ�rø�O^\(����.mY����* 8@���?\ ˰bxCM�ю�҅@Ā��Zg!Qp�˥��%�|k��b���p��GBlu���*���cF@��}��N�I���	�o�V������{D~��m߻��7��l�Wg�_7N�:�G�Bp�Ua)�u ��~[�6J�~��0I8�П���B��)��X�p���{Y��ot��v(�rd����I������%�JbJ��LS��S��qR���㥜fy��7�LG83�qh5P������Y)�׹]蹧��A)�2��ۀ�Nmw��;���Y]�8oc&3�1�ؼ?���	ҺA�~
[~?�P�\����6�EO<p��߼~oR�ԁ����ݓ�wwh�^�j8^9��*���c$���l�M�՗�g�&^���=0E���L���bC(�V�y��q�^��ǹ�0���f���G�P&��Z�1�%���oݽY��1+O�ޙ�a�z��[q��˛&fC�u�PZ�� Z=�ɼϣ�aiw�C�q�2�ٿ��!����eb!��Zg�]Z�V�q��0`;�.���ʈN0�5�N��xq�S�LЗ)�о��b�L/��́���:P�Jy6r��vu}!)�A� �S%������D)a%�\,'�޵"�r�Omđ�0H�H��h���p+u�5����R. )On5n�&c��D5��P�Ri0 ���k.B;�v���B��JD���7z��I\���Æ�0���H��U���1�zkө�E�E6k*x�������{~�=e����Ѫ���B��/����$в� 1~�B�=﬿�}Mg�DUU��-�J���0h�Xq�����t��������M1f2�@�[�Y&j�`QUP�A�taO�ɟ?v23����������o�4��S�,�{��8���-���7�*0�{.7X��V���h�E!{eVL ����P��T�B�*�+g|�t���rD�(~"�q�M�l�mHx ]�n\wngc���R4c"qf�Z������3�I�yX��_�v�9����9��=�V�B�X_���'�{�%e����=��_>,gյEJ-�N�WtFIN�����#ܘ�k̢�35b�aQKC��ui�+E@��/(]�n��3x����gs#���{6U8���'RI<��+H)����L�����0'�����E?вF���X+hu�p~�"Kj�fډ}f���NyW��\v�J� ���J:�;�;8����:���u�I����P5���\�k�W�6�X����!1�Y� ��2�ubT����n�����h��ں�Ϊ�S� �1 �H�����_�_�u6��	8H�~�f�d���Tw���C(�bay�ͬ�1v�0��|Yڞ�#a0�nR�;֘o<�b��~�#d�?1��giXR�[���"Uw	��̔�0r��U,�ܽv��М����)��.	�s>W�"���0J���K�B	�ώ����@�<��F,��褶䊥�!_By�õW���4��w��*�[v�����K���{�P����=F޷�����ۜ������8De�����m�B���{�$�(�50�S~b�4hR��o\kY����F�r9��]DM(�[�3��A>���QЮ��7�j�z��t���n�g�'�R�^��(�n�w�� |\V3sX�&hNs������X�	��7Q��1��*�\�VM!.�F���hMQ�����9���;pm���  �uP������n�W6�,�N�cZ5�<���y�5"�`���#�x��:Q͍:S��?�{oO�(O�_���	BR(F��nG�����k(d1��nBx�����#J�󌯹�A=��f�!Q�e�Tuč�\�C�@���|eWs,m��~�OF"]�#똸%��Bk�x���X� +�t�N��-�.�,�5����g��X��,��rB(uF��e��~�����\���j�Q ��^��b�=����/��؅���Ɩ"%�	�����E�$gNwN���>s�TQ�+���e�?��֯�p`���C����?&F��!w�.B��Ki�͖�M�Q�6��	�ؤ=���(F�c3��xu����b��ȟ����fFC�t�Hj��X�5fׁx���L�
N��t�ک2�뽑�n[+�Y�gQ]����YG}>���XjE�*�؂�Q���*Ԇ����#0�;}���I���鸈q����A�_��o�̟�G���rw���8dTՃ�s��R&Cc���wfK��q�>�J�H�5F��r��u�{�i��译I>�~ Flb���L

�Jix�!#�`
��_B��h�v�F�bؗ��zv،\,�P�/2q��w���Ό���X�z=��3.ᕄF�����P�
(M�/)�9A���Ͱ���}O�=j�6�H��p����x�!Z+��[����b]I����z1�}��Qp�'�z
}'�q�y������j*{����� �4�0�y��D7�K��Ϫ�":��;�`@�e+a��`�䦲E��Ɠ%ʬ���z/"�"ڍD�4�o�
lXko�e�Fȳ�-a�P�@��ɐZ|�'�mW}[9fH|R���,^��-�c�c���٧��aHŹ�ޒ�k�[B�������n#�9�zf~Aܹ^�KM�ܷ��W��zV�<pE��u"r�
�
3B|��ЭiŎ�/HB��UCAݩ�ؚz���ņ�X
_Zt̂���ѢNy�ƅ챀]��0����%���R�Y�Xdj�\m�̂�dO�ɲ�-
�<2X�KWR������+䫁?�czN�j�+̹	�i&)�iVRn!�e�s(����Z���</�I	CrWC­f=�����5^"g�L<��J�6F��~����m�_���&Q�q,�h;�*@���,�F�O�'���	�Xm��v,D�ѪÁ�Ǽ(C�R��~e���T.:�)�z)M�h@,��Ȏր_��轏�ǈ����V��+�n̑�"OHjDfeɝ�����t�<�3��Y�F-G���R�
�+A=���԰vȼ�[��g-�t�aWvH��P��,�É���n[��ZAm��K3�kK���.��)��w#���n�<�qE;u	4}�'b�>�_gp���d��Ͽ��4�üA\��ՅCGn>�A�َ�D����� |�I1rE�,Qh-��.�	�Ø����s*D��,aY�����t?ʷ�t�f5�����8��or#+oP�2�J��¹��JM����ja�)z��8�J���WT=����#��1>�
R
^}f�������'����WB�9��2g��*^� �a撱JgI�FM��k�"RQ��n�u��P�>0��;~�{�9H����!�]�ϣ/d�B��
�GL��.u�� �c�O#�����p?�oۡid8Z�6�v? h�v.N~�z���og-U��kz��}X��E�Ё�`�2�1��2UP�ֈ/�	�ݲ���xw���d8�S�߻�=c��gu�Oo�2���U���*�a�r^�������oVd�4�p� 6�{w�&��h������=�W4%��*�$��؊5�S#D��ofi&
�W,(2\�$Z��C�@C�����Q����/���hV���y�Y~揮L<BW��1��U ��@�PfK��%��eUp3�45)��#��P\`Ծ1���d�^����Q�� Fb`���ƥ��U�:ow�G�D���k��c.��Ra�\�ȱ��ey ���0lq�#���K��x��sX>,n���Ȉ�=|�p_/ꠔ�[:�1$�@H:��+�8���xG`�'{��SX���"�Fѵ