XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� T`}�bCh�J�������=ɀ
EJ��l�)���Kl���_����Ч��2�gg���L0����:QI,��z/�3��"�l��,Y���V"���O��L��G�}i��	f�����*~�,䄦�1�+.�̸ fX���u�:s���A刨�u=�'��@V�� �y�X �>o�����>Y�yS���ލSգ%��hĢ4D��Wgc�u2�<�� ������b��0c��<�.BRL��i'���%�;{����k�-o
�c���T�������6�2yX�����fU�x����8F$���6�|�ҹZ&X��/[LnQ�����$k�>�p�T��+�����/V�L]������y���2-����ɚ�kF?�'��8��y�#�fI2T��5�C���Y&�5A�o���<Jh'�T�t��uUM>���҆��IQ��P�g�2sũM9�;�C�BtQ`8�=�ŭe�>*��~�K.X��t˃@	`���<��q�?�}�C^��i]ٿg-t�q���c��1����E�ާ{���b��I���`)B� �jkN�����a&��|�h�6U,_0�~}HU��d���+��)v�c�����E��ΫF��L�E}ЈI�D�.~�Š�Q�c�s���!zz�c�,Y�v�
RJ@9*&��^�ϙ}��y�,"3Y�2�ߝ����;�(+�^N7�M��49����A\���*�4�D3q��!�h�z�˜�9�Q���$�6Q�`+7}@x���R�W���XlxVHYEB    3e51     a10R��	rU��h������΅�qK(Q����������cp�-�?���y�����f8�ϫ#���Q��": �U���S|���:;͝)��b=����5|��+�3�j�̇3�����l/y]>s(���s	�R�`P�E�kRF��z0IA����wf�]����y�!���[�t2c�'�e��_V�)��z.�vE�x�_�.��J�`	�,����r�����z���Ԁ��Q������r:�J_5Ș>֊c�YJ���zr_j
a�C&�sS�e.8ڱO\nZtY&���{	���*�<��1�(?O]��P5��s��Jܝ�CH���T�K��o��U�9��ˢ��{�n�u>�?|���Υ	W��7�e�\ ��-JN3g	wwVMUv�s�5�7�幪� 2wO�D�ٍ
�^�7��]�I����A	���0lX肞[�{}o��?�	7�M��8cQ-_�i��4���.NdBOy��&\�-�>��ŤH1ک���4�	��bԗENή�w@��T��e����G�٩k�\���J*���{ˣ'Â`z>��sF�y߸G�bDPC]�Gs)�0�^� �ԃ�s�p�HV=�,�f�6崼�?�����IJ� �z�j�';R���F"s�#ф���n�GN^*T��5��Q" ?$�ϴ�[���'M�_��/j�;�9ރ��,Y�цW)��5u� �vp���`���d��1P���X�V���O�	�Dld-��fӬ�,���*� ���P�D68�ˠ:U�H<^c�i�C��S>J��|����l7��OnX�����Q�Ќ��g_Y�(`��
o����ęMrP6MW���0�+�VlL�jSX��݀����S�:�y���&�WՒ���>�z�Ǵ�S+W,�c57�������5�K���|���[ L�Zմ/�Wz6�[\���Y�L�>�s&��ZT�T|�T�<���./?m�OU�����j�68b^%�I�.\�����X�|�S�����>�Z��VR����x��^�*GR �EսE1m�̹�!���}�Z6��o�Tx��b����D���.~8�R􃟵к�P�sk�J����I��H7/;gE(���2�X���Wl�h#ê[�ҽ���;И�%� �~�p(r�r�q��Q�چE�=�s��[Hw��?�k��±�����~(���a)�����%px?tLeR�����L@���}��� .O�^��X���ȓ�qSBX��*j��O��n�u#���|ش �з�m%A�G<8,]����Xou�@/��Fbf�j!A�<:J���7][ҎP(��+�Ś
EcMG\�<d�9�to,)Ͼ� �H��ضoΖ��i��������	N�s,� 0^>3`�Å#�b�:V)� j}�jnޤ2Q,L����5�ޖIz�9k��վ&\�E 7���P�`�	>���ZqOo�̒�O�v��|�8^x26i�OR��32�N���N��i�hZ������&`��?`��Z&����'+c��JmCS�,b��b�h���L����J����v]:T�S,,��,:�6�'$��_A
��NGC���w7H%�y���-B0����[� ���Uqsz��D=o��0Vn` C>�U�y�H���B��>��`KĂ���~~��ck41y�Q�P�d%�I�vV�k�t]R${LW�:V�mF�g}�+Mol��JC*�=�nW���$�s��e��u�Wהd���}�һ�9�`�e^���傽��:����t�T�����sD��comhAe�����H�?�IZ}FsMӥeȠAț�=���l�Շ����J¸�<�r�?�>rl��LGC�E>N�g�����jG�~�2�:��,
���˚d-���}�oV������*0h��-BV;�M�xR|�������͔��R�i��t����e����L���>��<�UAH�S���-D9o�� zo��e:��~�"���4�B��s�&Ӈ�#qk�d�H�c�_��%��P�Q� �Z����,9�.,{�`�	(av�`Ĉ�;뚶��q��Zx2zIb�YmtJjm%���W��&g�gv��P�!��&�������5�A�³,`��&r\T:��z�v$�LX�����΁^LH��Ћ���O����8??h��/ò�v����ĉ�E|�E�/ԦU�č���Lݲ��o0�B��*PX��١�M;̐D;h����6���o5*�T��{qe�:��<'�Uu���`iu��^�u�0{ݲT���D�D �x��+���ß�{��=��c'��q���g���i�-{^����Ϥ�����i�1�n4VD��z��D�я�mӇC�"� e�M�1a-/>���]�1�OK74鱗.��aޟ����5j������Y�Ck�T��4B���!��v��٪��L�/��)�>2��3�w���xH�Tf���tl��t�/P{�Bs�w`���MÀԉ |��҂�@ݺ����_¬�����H�