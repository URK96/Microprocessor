XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� +��@Ȃ��o�Z�1�\�s�Y/9�J�æ��X�╚�xf4[-A�M	i
��,�d\�^n_7�Ⳕ�2��~w���ݗu��j�0 ��,�{(1(&O�^P�u�\��^)I�%\~qYS'^0ϵ��"������y�J�rg�0Lz߻�Bx$��d;�]JJs0����K��/������[c��mL���gf�.��z�w��	���n�7�i��˂�>�����Ч��{ޞ¾zo=�z�M1W9��8sNW��NƩ����s��4#/pr�'Gp�����/���
�f��g��bW���a�Jg|�|s���,������,J'E��lQW��j-��3wR
��/����\����(�bM<d����X| �+6,�����qgV;G��[Ssmc����g���B8̺^��)����mNݓzBDT�lgª/b����2�V���n\���^	3Qq��z�WJF�B��G�.����Z�j�[{�Ԍ,h{�'3�R����y�;�9�����8D�/����١%�z�u��x��"]�yR�v���+(NWۥF𐡷��>̝��H�b��0����nk�5�`����HD��RmV��V�!k����oY�� ��h���r�$���&|�O�V������>��ڬlW�-v�]�%�UP��3��"�.�����P�^˄� e&RC$� ��K�-��u�+8�.��=Q	�GR�5𴶓�����Y����/��l��XlxVHYEB     a56     380az�ʆ?�c�&ڂl��8���u�;©+��a��&F�5�;�����X��aU`��w�at�s��,Ѹ<7��H�^g.˺�ԵqV�����N?{�B?��򾡒��c��_�8/��|�
\�g٘-�U�6�+��U���8��Vy�1'��Be�7`u��[��1�y64�Ms��C�{p��'˳,��@���bE<L��"2lg-�)A�qu�1�V%2�_�U)z%d�\y�>N�N��~wxs���Gb(jd3�UP>P�-;���T`&w� m.N	� ��a��Jr`�5���j���R���9*�Z��_�C):�k����N�	�w�������C���<v�
Oc�>��*�w"(_�"�W՟+l����1vJ�˼�^Ìdj�;��j%jè\��2;�����"k��
�sXoF����������az��s4鞁��GU\��equ1ľf#5��ɶ%W�Tmh��?R=R��O�W�����nxQj�
D�)0Vk�X�A5i�V�� ���6\��}D����5~08�"H�s�I��q�l)[��$��n�F�	�Y8�E�Q�n:s�w�	�N�\�E���n��\�-3cFe��I&��{���$�f\p?(Z;�x)��tX�>c��LaS�5'��k3�]Kٶ�ܞ��T��ڸ+p9�V��r���E��/&lV0Ag+m��t.�h�����ח�u���>�m�t��-��M�ah�� @��X;�awl�-�WN�g��t��ߴ@�r�r
ʣr5X^b>��}��dN
��a4���L \��r�ч��l�c���T'f������Z����EK�K��qJ�,���䣄"�4Ɗ�S�b3+�~��b�����q\�fs�i��HH NU�������Ś���-