XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����T��m��OH:!9�Nhg��O���H�WiT>��{��+����W�ޗ��v=����g� {�t[Q�0�Β>�ں_���+C����q��1Ƀӭmi"�n;���HQ�u�'�A�6���L�Mn���I����Z�#X(��Oz�x<�;����|Czn��"$���`�}$�1՚.�JT�v���x
�0 7�r�d�ԛ���7�σܝQ˽�4���W����E��^hڈD�G��v?�W�S�'� K�O�G����������ZGfk�W����|T�����Z2��h_���?�p\��{Y��Y� z�Wh���������O�FK�owINU6�n�3���h@yJ��&�3s{�g7tb��0m_�Gt�w�j��eO���`J�)s[�Ȍ�ڏ��_��g�"׼mj����G% y�M'&.b�T���Ķ�*V����%�G�� ��f�����#��lb�m�'7���Y����c��>�
|f)�XsB�!�M@"[��jؔLGe�l��5�Y`4Uf�~/&�N����wi�Ny���3�޿Fh�A<°�H9�i#���׺c��=��NV�����;Oz�]�=��x��Nr�鄏M /6^�
��Ŧ�0�"Z0�=I��+l�D+�=���p Q����cᓹ)/��:y��ڈԏ�.������ƴ�P�b�p}'(�پ��R���5��-,F�sC��e�,Hx
�ٗ�z�Ha���:a�����P	��:z�~���>���G��XlxVHYEB    1cf8     790nO�|d֮�/X��T�`�B����IE�RW_�^�$��>�V�a�"�n�� {�LV�P�6�(���.q7A$&J��>q�<�-E�9ƷA��x�TfHTM��I<56ioq�W%��٤���r!~v����9�ȞJ��뺃�ҪR�Fд�$n�� ߽��%�\;@٤y��ƬB��Ӌ���nRC���l�T� r���/�;#bTPC��n���ryւ��9�7
s���3�����a_j�t1�/��變�`�H���`��Aw7\3���ڡ��v�J�-i�XǞY�D0�r�&C7��G^g�Ⱥ��)�i��~�_D|��M�p-2Z⶗i�e��C&�Ykc�I{�"b^�C%Dz����'	�'Y�@'����3�(i{����0���1<�u����
�Q��eh�o��&⫶ Y���:��M�Njxv�1LF�8��ԑ�ݺZze
.���;sU�͓�Tj���Wd�b��W���������InQ�H��ښ�/���Ê�}:�W��Nyj��x�����b$)a�:���ޙTU�B$q��t|�<�+��i������g�1�$\��-#<b������(TH��c=1:1���Oj��Z��T�d���&Pz�C�h����j��D����I�t���1��e�WrþQ@`�-`�%گ��]�1����x��N���&JJ��^1	!��PY�. ܜ���=��D�,�zt�\��.����Ԥ�P��04E��J\q{`�����칉�գ+���r9W���T��ūT�XHod|�0Yx���pu�sfV�w�Z KY��.��v(�܁/���w�F���Wܑ�8�Ћ��M��
Xh_G������b�M��~�Lw�$>�F�\�q۳���gW�^+�d3H�k���_����(*��	�tWm��7>5u��é��|x7�k�ے �畉D�6��C��w�1�z�xh��@5���$5�oǬ+���0�]��s������D��&Jw=hGi���5��/�<����{�5�.�ؾ�ʯTz]�.,E��>a	��� ��V��m�gX�4�Z��5ڧ�;�����v'��n���ΰK�vBv��]#Z�2ڄ�Hg�yH�><�c>�)ط��ā��=��29��H(�K��\�ß}6y2헎�|t�����W8]�?h���CV������?�k*[�̈���V8��-C���ƅT�yI��cA��

��z����uт�;�9�FP.�](�>�mX<�>Q��'�a$�!�<R_�u�c�5��$Ħ3�Ud��"G�#��R�@q�Z�o���=p/����gU#t{Ν=��Nq��(�Ϡ��W��MT��J�6����*g��M�s:�����Ýs*J֬�/g�>���+�͎��N�P ���[b��c�S���a�-y��=!�od,Wk�Z7���9:�0�.?�?�%�}�D~<o��D#GH��XĬ����������>�fÈ��e��27�K�8P}���,��$�;N���ݻ%�Fc���ܤ7m����>cLBO����4�FZ���$�j(ǜ<�A����O�����l���okN�������KX�F�f|Ǉ� �v��WE�?t�:vh=(�����xd��G��YI���>z���B��E�F����bV9g�.]�Oh��%�f� ���|��V���ƕv�7[�-���=U��{;,ô:q
=�� ��J���u�Ld�Ͽ5	� �O
 �:U�B����y��֞p�ܮI�d��i"LΨ���u��S�b�!�4w�%���B�k1p�p~�������i3��8��>xτ�`�1oEdl�	08��5;]!;�7E�