XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q$�7�]ʠz=��.XeϱY q��;7�W���^�ۊc��
	whD�\ⓤ�:y��~�8�&�W�c$��>�c)Z�u'�(��.%����:��J)����s�G�iG�[D�3v�h���i}��~��߳�YYQn�r���a�n��;c9��.�Y6Ĕ�kWz��b�8[�?�jW�d^=��{�t�ӂ�0�R��~5l�=�vf{�p�5��/����V\hDO�;@`ha�=?���4�v>��"����r�l��L����E����,�u�!�����_�R��g9�x��J��b��=R.�l�+�Ox�h��aU?�-
��<�b��3�Fw_�+{P�<��a��e��[RYk�&�@����b��phȀ�&ۅ�f���~@�(���9y��d�I�5���Nh���, ����{c)���^MG�v~�ut��=���g��+�P�����%�r�������h��&�e2�:�7 ��і��).�n�adKn?P-ܚ�r����������L� 2IJ=g�f����<������3���Nu/*
�$�2�\�j��C�&����FJc봩$R���)��W�	�3n!���8��N����6uT�(��n�!s��3SZ��=�U'0p��"F�{�(�F2Pҏb�yz=c#ג��w�P-�W�;�]�B8�ɘR@��,{�����E�Z���U����H��l��a��{b�~Z
�^���	k� 3z ��/0� /�XlxVHYEB    1901     4504�� /���b����W�'g�T-�\��)eAB�hј�tE�������k�@p�����\_1-�p���|�j�6�}�`��N��lo��X���w�ow�z�K�����l
_IX�b��`h�ԌH��H�:��
( )f���S╠�6`�`-B:N{ކ���q_@�8a]4b������ȹ�!��T��P���Z ��0)K��@��$�9wv�@�W�L��VSѰ f�f�/p`�ݜ.q+���`3/���_S��d���!"^�:��OY�9���'0:]����:ٝjGL��L�p���y�&�"0����9�U����&�2�D�U����uh�-���}�ڙ;'�Q���<>Ɓ�:.qa$u�x�p����T��ɽw�2���I������Gp�]w���xhs*O v�b���ʞ� ��4�������O����/z8P�48�a9�_�*���������D8�IAz%���YE����@�?�]�L�����EE��S�,�f_s�ސo:�]&�O��Jl���	+�����zr�K<��bi��W'|����8�G�W߿��/��9e9�-m=˻2�Q�����._���������� �e ;��ѡz�Q�}?"��a"����J�:	Lх���X`��~!5�����2�:��
^���{q�RPPǔ��!��LGi+���X2O
����˫ͮ7 v3Vo(�VR"a
�t�R@,�6�emۅa�t�y�T$�Z��F��q���q���V���l�äȒ� �ς5�Ӳ�qZ��N�J\�b���nxZ�1��A��J/��x���ߢ�Y,��Bߦ��p�Z;� 
��ǡ����ǒG�0R�ɖ����K���x@@��IN�Z<��o��GC7�@c�"%���Nz-}MA((_T�0�i��d0.�3y3��7���설vj
�\�[]%�ʉ�Q�v��:U�G�܃��hj[���x1�怐�� Y��~�p�Od�H�e���kdBcnHvu! 7-m��-'J5�|���R��8R����xB�Xr<��@f���m��k&���)�����8���
"<��E�T6\��ӹnNJ4"=��