XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����/4�p��N���(�N��]@v}�N-QA�v&�X����|H
�
p�3�.E�Z��?�>o_Ä�����s���m4e�LF]���,����|hB՛B9�q�6�1���o.ec!{cy��Ϟ���fFȊM���{�U��D3�	6U�(r��1�ʝ�Rq'Ό�:%��C~ ��"Z�:�gV�=kq=-0�I��qA]��6�����N@�?��<Ƴ�
��i�UGDS�r�ٌ�����w��ψ�2g����!m&tS��ƍS]�5;���H숹��*G��Ŋ �J%�.�+��0��Ԙ��{�T�J!�m#��dK�ޟ!��1���9�@ãp�/�Y"o����и�m�mzXT�|b�G��B���~�,ls�����7�O�\{��ɬB�Ѝ�[�ZG���8;I�L�Tх}b(�x���CS��Ӑ_��v�wv^>(�˺5�~��Q�=T�0�K�;���(� t'1sM+��6�+�F���X;M2�dC�>���#~�:�h*�E��F�[��$15>�QtI���sl�jKњ9���'.G��]���
���t��+�T�E�l{���=i�G�X�� �I�jQ�UB��-�㶨�<�� � �%�>�4b^꒡~��1�2���|Rzz"���A�.c�	��2r�1ҿD ���9b^r�	 ��`�$ѿ��q+*�J��ۏSe�[�R:��l�ChPܞ|�V�mm���f5����e��}�(R��bXlxVHYEB    fa00    19d0��ķ����p�\r:,~���eu�`Gt�0��)��r+���3�4�h%�V.x�GAܾ����<u�����&.�|�Ο�7�' �k�t��@o���o`tޅȽ Ƣ�!�9\��nȕ�i~>0�T��e��x=�����\�:O������+[�uW�C���ϋ�,! �#�߅1癄����"\lX����#\A6*��R:��nVr�z��Ij~ƞ�;V&��}�K3��x�� ��o���sk�]�\��6��e_q�H��V8�/���R����f��ے�s���;!���[y| ����K��_���TI���nC	��6z�&�l)M������i݆=��E@?}[<n�辱��ذ*1��mXM�c��@�}�J����z�G��v��D�Y[�t�"��g�D]g�Ӣ�-��G;�A��0_�]���.���{��ϴL��0����s�O@������Hc�.I��8oi�%?����JڌX@��F�=�Q�Xdw�9i���	Y0WԺ#�%�@ �?ʹ�YW�8�̓P��^lY�;TG����ً�^���_7r��$����Ы[7�9���>��W�a�8�y�C������2BU��$%Ł��|[�0s=�L���֬�q�fpV�/���F;��r�C�ͣ%���c� �^��i?�ا�d1ܫ�
n���}���#u�������cAJb2 <_�,��7̾=�{�ǣU��ita�*��״f����1�n���N�c6rV`=������d�������^! �����;1�"���	���S� �cגf�����Q(	R������K����6�q�.z�f3"L!���n%�
W|�����z�	_x�]������4����s�sEf��p�<&*V��?�_��G
����-ބ�3=�������H���}��=����e�VT��fЍ/'b��<�70 �/@�a�	iԦ�3+�ۜy��q���'�oUR�0c� ��I[H-E�,MQ$|]}2X�u���·����N�(�"�D�Ŷk�h5�'�`�,5S�G�wmu��ݳf[�^zK�A��,�3�dw: �S����*K/y$�������
�D�\� �a��0��7|���V����J�b:	X���*� (�o���k�0��w,�B]u�s�� � A�K�1̱sq�Q�[æV
)9��۶�nt��ҡ0d����L�γ���Ss�5�)К/���q2[/�9z��x��S({�>d94�iI)����RX�3#jțWz�薁!�I����?�6����~H�|�'��60H�b`~׊��3C���Ec� 4b���!~xy0>	EWĊ��e7F�L�)�X%J�����Պ�kp._��YT��N�Uc�h�g��4�G���;�!����2}ҙ07�p+&�m�\��ݽ�}zm��ZZN��@L�۾O>�rP&'��s�_���6H`�4� �.�����W1��`4���a(�߆Q���׫igg|b�����˘��1X c���
�g�L��/�9=���dQd�|�B}����o�Y��l�#���l#e��k�Zq��>�7�yq�/����P�p�]���@��?v��"��T}uQ܀B�/F�%<�%3
5F����#���ʷQ���z�}��ہ�s��8�b������p�f}G`�\/�qj�s�¸�T�ù(�@*T���L��aC����7��Ι�0a��Ԉ���M��"��:��-g�NE�����̵C�}Q5t��!)#yi��R�[e������p��v�pX�C�P>��ڬKǀ;�����SI(mvxu��Jv�U�s$�t�'�?�!!�Ю��d�э�no�GE\Nݩb��&P��ԿT�I�/�'�f�f��������KHJ���{qmh��(�c���~un�_�*f'�O����+���҉�U����Ԯ�����:��Q��]�]��^xQ�­W�I_VA�3���n7ՙ�~d$�l?a�FP��%���R���F=(s����}ٍ���<ll��n#W�S�3��@qj�lLDn1U�R菽���6�&B����oq�n���0{�N�eO����V<pG��'�Sz4Ox'���r�f˷���u�6�.ԭ%��kx<����J~#{)�����.V/�$�x$�;�t��L�&s���yKհ�2�0�{�x���R�����]��f�ߎDr*���h��ȷ��@@�Fc"tZm�,Ҙ%�h?�F�^���� ���D���'6X�avx��8��;#Ke��g����p^F��ޥ@4���+����̥��Q:){`�=) J�]�䵨�6�*3�.g��Gm^9C�O����ہZ�0�������绵��s�a�%�v�Ůd��m��+�T�{��\�x�0�5��|=��rY����P�
���Ki�S��Wѐ�6C��8_&B�5kt��6ʹ�wC�B����駕�ᜠ��I�i�� ٴe@�uP�!x�5�D���� ����B�?��a� i`T)�z�q�����v~ߦ�����>��W��"q�2���`�$��v�N�ZaL�[ hp[���T�����g���k�l�Cԥ���a�Х���*j'SjiU#�T��*&.Lt�V8���	Ȩ3��֙n����zW`b���dx�n6) �ë1�
9`n�z�Y�.%��U�)�.T�'�e6 R�z��g��$;�E���R�ۣ�A��$s��40\�� �Ɵ�Rc���YH:��lRG1�G���3Z5�V������g{dƿ>s��ԘE2k�f����گ�c���?[�{o���� ����XN�$� �4W3� ��4RӤ���Cc%~��1Mq5�ބ�����|���	�V���z�Ic�>��5�䪻����%X��=`Ў�������BZ�5�0��e�����ݯ�yh�z�	0�8�'[�(i��'�d�h�I\0zHfZ�%�63!	��5[E���b$��<'��i(�f�#�!M��;uJ<T�6�D�N�dSW[����ڋ�x�!�����3YF������Zy���Փ�HGl䣝����3y��튣��[ρ�2����v�ݿ� ���P�k�-s�<��_L\{U�j{2pF��PӐ]���{��^<����և?6�J�'Oڍ_����$�Ej3����`����b��V5�uf�����f��d�P������n0����-�M��(���bS��M,�_/�)*�ؐ�?dz�=�I-� �i�7*ǅc��)\}�Xyl{1�9{��Ґ�\Ϭ�ڤA�1<��]v�~��M/q�h��Y�*��EP���~!�IM�~ C�Tm&�:{��t!�-W΀���Ѐ���|E�� )�ړ��ew����xu�Pq�,�u���|�I'�;���Di/Tv��4���A��z�5(�c@
sy\��i��5���z�Yc�6��6��W�M�c�j���`�.<#��w�/�D&?��m�o�#���r� � ��.`j�}�� ��h`�銷��S.��ϔ]#(T��4����ƬB�zG-��/p�E�Y�t��fW{�v@w7"x[�C�6M��3Ț�A�rt:1�-#��o��>/n�wŶ{�g(D�ȓ� P���4Ę"�T z�f�6`+1�a:u�Tƣ���F���*�*��]oD���^��h�W�Ҵ��z��?F��<~�k�'Mo��B�7_����~#������^�P��k����`������=Hgk��_�<�,zuZ����Je�r��7�?a)l2��|��'�/^�;�9�����h�dgd���{�x��A�/�뮤$�;v�L�� wa��{�G�9�������"1��"�֖i��|-���(6�"`*[F�V�%��D���h�-h�]Ѭ\:-�L�6��l1���峮V�&��Nc��3�J����ߜ�(�����$�<%�r���Φg$�X�V�-� �fZ &��-#��C=<Q�g�f�����XPOT۶��r�LL��y��R�D����R�" D��X��Ar)4�����6�o]X6óW��.��Z#,�4�@���#��Q��`����5x��Q��	�6�z�iX��c���L�3��~_���Cȏ�9������>YS�9C北�nH<��~ fN뿣+�TZ��@�P�����y�������>�ڏ4R����n��b�^s(D��iS���{O���e��X,,h�62��.�Z�j6�uŊ!��oJQn��]�9�{!K��;�,�3H\Lt��F��[�Ș(>4m��k�������e�Ug&�+*]a�������ؖ�ߕ`�.$YYUAi��y��u�ȭ�m��Ō.�6H���f�	��E6��8��3Rw��t�<
�����J��'��>5�&H��n�"�^�2/[9�A���Ջ���������X'���!��Z�1�<�
�V6Xߠ��JǊ�
�$�v9�����	�u+���|�#�&�&�lmO4g{y�qi���>��k9�G��N#%sx�zpz�Чdv.��a7$���A��0��誻>�A�ER(e%5�:8�����$n9K���X�}
$�t����O��	+$?C�Ỽ�x�W���6��[� ��r�=��_��Ï�;�y+?�H;�w��Id䈚9�|h�i�I���zQ��TNB���AES�>^�%�+��L�Q���x��l������+Ҙ�ߣЛϾ�Y\ �hq�P5��I#�l!��jl4is�⪳��O˸&�!�"��܊��KO��ܯ�9�
��M�)��9D�jҙ��=�S���b�aH�Qcb������-J�*a��a�� � 
��d~[W�� ����q�g���t0��BrYahv8���"�IȠWOϳ�q��Ϗ�6�S�"�9�KV��$��v�ȭ����r��L>���E��3�V���!��\�(+
�<HF�6�`�6�7�CC�������[�������:�L�ý܋|�� ����S���#�1�c���t�~��Z>���QV�}M"�.d/m�F��/K��ѱ�%\����[���B���q3B��=�6�+ƾY4~�>��:�Ɣ��@O�@�ė]
L��J-��X�Χ~��f��}��uR}P����|2�#Τ!'w�pvV�
W�hzY�j��]�A��B��[)[�f�7h7���4�4�e��.�u{��򨅣����P|���3�'���16�\ ��j�u��x�?77���
��v=����(�R;�v��ߡL`6EsMǴ���
�����?��u}����sKJ�a>E�_nѝ�g(���@�!��e�]zb�Ǆ�n�mU������^<��L��x�ca�	�	�C�dF��f���K�/�.�mE.�K��w�n�@+ūtk&�?т�V��tn�$�Q��*��8���
p<�����xTx�Z6���b�����ֲe�Q6t�X��гA�K'J3�f��N��S�I5S�����8�f�9�t�nE�� h�M�@H�����g�.8f���~�=��G�x���M ��3�(Z�)��=���P��nUyU2p:d�5���L��r˽jK񺝱�d�1>�-#3,>K���ё����g����5�G���8jz����؎^a+���3�G��6a�-��`�o��E&��mz9�{�����j{j*�ӡ+6D�ٰgK��.����aHQ:*Դ���,�m;��g�N����� ��H��lb��#!��{z�Ӭ��S�i�/��YN��
�)���u$ZpsilQ!�*�c�Z'n��1 Z��3/��ђ�`�����I�[|'c{9j�iK��İZ��u�C��%�7v�y�����8'ͺc��\>����A ��A7�X�Ԉ�KS_��YU�(�2-�J�W��4��.$����H�Po7�P�A�q����C���sYU� �w*���P�
u�l�Ǣ�g��T-l
"hބ���_����%��(|_��qiU�'��z��%�k�D�-�Q�\�D��/���t�'��țg����*�7��ұ�E{`�qO5`�����<jN����X���,֣���-T�M��I�}���thZ�Y�E�upR+[h�D�Eۉ�u_��# y�BP�4O[X2�(̣�'o�׹��]0D[�ט+,���rK�c�3l�.��Э 5���ԍ�|�Q�?هƂ� ��*v�d������ 'Aߏ���ńO�뙓�➪d�#�O��6�G�������T@��n�5�L�Ƚ;tn��?�A�j+��Vv�Q0.�6{Ij��������p��@��W�t�D�y�]�t)�W�8���T�����ޕ�N�t�}��\N��N� oa,�Y�謁�K˂c�����R#��*��%�J�I@ҥX������1~XlxVHYEB    fa00    1630���ORq�u�����$K瘣WdT�4\�l[%z7��2������z�B���]k_��iYP�9g8������/��G�R��+_�1�ѱw��3�醈���<�e�f��s��"��o�ؙ�����96�HWr	���>d���۶F���"��S�;X
5.��=O�7��Ɋ���Ф�mj����!����,z6Gm]�$l�4� �� �	,ݢK�j��h$Zj�a@Ĳ�������	��
���x�?����-#,<rx��d"Dc�}1(k�N�F~�+��\�8�%�8�Yë.-���I�u�z�˵y���f&7���NT�{e�ǲ[��;��ºú��:%��.��#R8��T�U�>x�/�}�����蹇�v��äξ:8JM���N�t>q�<q$ Wv3;�,���c��}i� ��'�P���Rǁ�v$�(��`E=�y,�����n˝U���+�v7���:yL��s�yK��r^N�E/q�Dϕ�*���G���x�-iY/�ϥH5����͌�}UU,J!����![�!h�(����|tp��T���3�����ήU/��|[�n�O �t����-�*2cN�S;��]0�s����� Ƀ���X�ϥ-	Q{��)D��[ۂ�vT&6�}2��O��2_�;>��&R2�؇���ɀ��d��\?KL��Hu�[�m}D����M�."S�O8�s�r�{F	NU��Ų�/����ro�=.�'$y�nf�xBA��PdT�ˀ�Z��~���5�7���Ys2���;Lt��+/��^;����3w_�舡�s3,J���w�JK�ly?�c���{�ԧ�,���^��J���7SXʉ�p'�/�m}K[~siS�I󍨃�y���Q��A�,i����˝P|�i���Ys� $V�R��`Lݛ�}\�xo�~���^uWp�;f{MB���0�28���UL`�+����������z�Uz�~�x�W��������_^�$�ėw�zZ��u�R�#�'^O�'�S�Z�4W_��)��s�2uU��Utp$ha�of!��:��"�����W�%$N����$5�<�O+�aι`��~YwG���Hl)�fv*�U<�Z�aj4D)�1~r���'bbg��Dq�[�=�`qDy�d�cG	i��1|�~�}H��M���1�8P�Ɛ@|}Q��ry6\i� 4�$�+��.�E!W���+iG}�׆F�qG�\T�
ox޹fM�׫���Vtu]����#���*Α��V	��x����]���y�a����T+�{�T9����_
��wHZ��Ya䩄�<��ɦU�i��l�@ %���4 �d��w�v&MXcWoXr��L_�ⒸZ��0�&K)�eB����;�M�	7���7��o�n�	}���n�t3��o@M�[�[i���&��vdNn�M\�Uǅ*������s�{d���w>�}��	�ś^_���⪮��;��B�s�9ȑ{���&�PrQ9T�,�P�+�[R�q�k�����C�4y�N�M�H�u{�Ӗʓ�����j�3ďg���S��q��0�$�6/%���Ǩ'LH2�ļ�5���QՏ�Vpɖ�I1��w�ޗ��u�k6	�� D�^}��*Lbz{'86с۬�b
����C��H��.Gvɲ�\�a�RaȾ���,�E����!��R�d�z=���Wnx��x�
���%P�#��7Y��6s�Dtv��D̆C�G� ̫Ms�s�7��d3Tc|㢞s�f���u%������ ~(>o$��<�g ��
�'l7+7G��M_eeĥGZ�PmM܇�Q�z��us�6j��:����o͘�+}ܓ?>�P ��*r`;o&�.��3�L�r�o 4�bI���h2���]�PgnK�?���h����d�z.&SNZ	�����?�4���!��rBb]��4��.�i���-"؂�9�@�R)n@��2iB�0�I�;u��
��7��X��f�~��C�r�	��d'��A���1,d���&����[�_%L�l���)Fs�����2�7θ�0D��"43�O��;1ɯ�m������)�f� ى,��6�	�a�)w�bY�R������b>;p��8qM�EmqM�QT�ح߾�i�Q'R�#m�� ���R@�Ddh�S]��uu,%؂NZHm��,�/O4�`ڦ��u�됻Bz\;UhE��t��	�O�	i��o't�6ܸJ�Z���U��i�fjj��9����e\�sU��ֹ{���(:�nE V#r*u1j���Z��K��ƙ�J�xQ8�Kș��6�>73�K��J�tì�äX����i�@��[�=6�#��[�|�rM�(K/
j1�/�o�lK�H�Mk�R���g���zxC#h�����.�D���Y�I��3�݅�(i2`�����_\�#T:D�P�b����_�J����fõ���G���Rl�5쫄UM�n���� �u�t������s��<�m��u?��B�	��G�D�1��鸴�/�Ą�n�<}��:�����n��&{���b7����,��"��<yoNv��L��d]�a�$Mb"G���t�p�e��^���1hy�	����	T���t��5�]����G��#��Pq�+�W
�G�n1������s�^�t�n��Ѡ�7���ֈ�i/ �[��❲��@�-�����_wVhd�EIo����gy9/���1L'�HZ�Ň��a�i�����8�<�ڔ���
���ץ�r����N.A��K��~q��p���fp��|+��7�g@ս�J�!G,,Yܗ��D_�]$UF<JnK�ialH�V�ܿr&����NM\�E�?�ܠ�M������B���N���8�xk�Zc�Vn�f�B���g���;ŧ���EJޢK�'�����S�*¥�-��LobQ���9Y���=�<^���Č��:����Þ���mXV�07��9D�H��6#��wn��~�R��7���/ �p��*��,�k��]���+���M	͟��w��2�#VPn`m���C~�ч^�|9�1��36l��������ӄ�>��@sgL6L���2���W}�,&d�&�)��t^�u]�v�S^Y��U�O:~���2�!Y�|����Ԋ��8Pj���k�\ٷ�xe���َ]31�wI�뢁莮��B�1�e4�XV:���x���U.b^��mݵ2lm�6���b!�~\Т�>Wљ;݈C��KP����}�uj�b�t�:���c�pr���s�!9��ͼ��0y�W�`��vMc�3�ՍQ�ĎJ{�A�~�RH�B��yjٞ���v-�M������p�T\J��=�crq�D$�0<2�5�:�����`�O�����{X�����D�X�P�4L���^*�&�{��s�J�S8o��Ǩ}#ăU�EW~�P\���)��W LI�T��s�<��.�J�f1��pt�K��i̢%����i�a�*­-t������{��b�=�rnD%�j/�#�z
e�f��QH�q�������%��D��k��fN��4�d���P�g���8fΫ�᳝�> wzL�}���|�G7+��̮�Ys�t;?�H6�:(���܊�KD��7����X(�>]�:s3u)�1`��;��:'/o�x3<��D'��h#��c�3 -hf����=���9��:hT{����!�a�s�gA�=�ͷ���=����Yd���`��.�.s6AW����� 9�E���B���ڡ/0�MV�vx�*=|�ǆk�$�{�
wV�5�:�]a��~ۡ�C�*J�_?�7�.�!��#Jx6C�yLX�4�h��TE$N����@>*���	���)���PsX�����-1@�������J1�mDM�NRp����7RƎW�!�gq�IP��*�	�Rg�#�)^�ݍ�Le�|�Z�ʣSxEe��	9����]rc�aN��>�GI�\u#�2�� C,̗���GWhM$�}HMcv�f�.Ў�Q�g�n9M<_���f����dɢփ� &E~�3�ze��6+�6T9��6���U����l�c���kT��F^>�/�ū��&��t��e��5���,��z�TJ�U�EU[���7J�.2t)HA�����:F�� }r [�l�kMGO��"3�+ǭ���P`8ױ2Ӆ:7�bs�B5~7�֓�Hc9����]��Je��ǌ����oB'��b����Ԍ�>�,�+A���y~���餚��%��-x_&���v��7� bmFW%a��i��"��1��XpWW�#��J!3������?7���%k����ScL�xk�l�D�
�+p:���I`ƽ��I� �l#��;5S}��K�:�&g��8���(O�M�Jp�:#�ej �u��y�C���v
���H��ތe9<-C4�c~1^�g�x���e����7��S�o��e>�G8��ͣGk�X�C���L��༚°�9q̱�o��D�e�e��n�G�6��|w��$��Z�oC��'�G�IYq��IP�Q�&1� �ڗ}	]�eȶ�v�*~>4*[D�m�_]4�T�uo���ʳ���I�%l�쑪 ���
���b*S3�}��{�u�u�	��N_q�Ю#�	����:����	V�veY�x�p)�L`��mw���Zq�J���mX��i鸷�Z��B�k���:K|�k��(7Rỷ�9�ʼAԜ~()�0��N$C��Ȫ�_5J^58;�ۋp))Cn�q�(vι�>:ɶE�B�R-�ՓN�%������}d�w��|�{X���0��,��$)�.�P~���V���9���0v�.����4�o�ݸ�0^f�i��v� �Q����5���!XCːi�*���]��hb��Zq�Z�&���4
�F0jYu�?��D���Xv[���?�F�&�#4bkl<"'0�6+�CP��r	/�Yo�#r�3G�[��M �5����b��F��VO@$�0��{>�7F醐�������$Q>�����Kh������\=���q`��}�0�'���0�2�JS�{gy�K����y+g�"����K�|Ōg�e���y�V�6h�k��G��*^�qu]&��EW�P�;_p�]�C�=sG��P[i����@��r�u�-U��W���	;J���bex��ǅ��\&�	��Q�/$ه��E�tpB	��m(J+w�:8T�۲N�[��j|�E��ȤP���B�t�LH���O|z��"C(i�����,J�k��1���R���h1��ʒ\�@Ϯ�I��o�	sM�#�HLREzV�0W(N�	��*]��3J��/U��7�ཤVD8�N��,���f���n.��)⬿�Py���6�x�����݌�r�pn���2��<��&�������� ��e��D��|����$՝2q~P�$�Y�Wo��Y'G�I罖ƃ���"�!��:l�</L�;����Ni��'7��� ��Te�"�}��9��h�Ȕ���3�xɺ������ԣ{Xb�XlxVHYEB    fa00    16a0�U� +8��R���~BC�/��qi#�u؇B�F�ʨ����+��Ǡ���F���w��Hi8��$ԻV��U�,�J����{.�_�d��Ъ�~H�Uҫ����upNڱ���OWg:�@lon�Z�y�K$�J �k�J��(�1�5�f5�jy�����I&��Z�TK��R�I�A]�z޼�P�+����̮�GO1յ9-�ta.Ǭ4��dX�h2DB��g2>?-�{�[�O-Ĕ������[�DJE��\�_��lf� L#C�S����|q�@Q��1�ޮ����6�	bh�2�X�Iw���=�$���&����ۂ�С���g`�,�\[�y�[�m8Ž���p*3�3Or�t����b�H��E����ı���Ny��ԹXP\/��'�\T�R�^r?>��kt �A��%#��� ӏ]x�j���<�su�� Z�F3ğ.����$0yp�=B&�*9�j����9>����P?��ؿ�MYP`��IP�t4��T��	Έ�40�J:%����`��>U(�`���w�N4UP>Z엨lےQ�<��KM�oܛxʖGg�9ةlV9�K.؈2H�Y�|�~�	m��Ww�ɽZl��6�Zx��U�=&��I�.�ƞ�b���^��xJ��p��ӟa ��e�qCh~5��3�<?�^�+����&�������a�Lv ��fQdQ��.>���K�ȻO��qH0�c���&�j�%��-M�<���w���dtNF@��,��۴x}zi��P�Y�?��E�R�rPM��#I�.Q误oO��W��M7���WZ��U��s��6�E&>�{L&�pY��O�)�`N�I�J���S�랊���9�\
��'޼/��@��� kA����h�T�� �i��b ����o��)���_����@��n'C�Zr�A�f�:���Ұ�����t�`ņ����E��5W�a���;�&�r��}QC7��g�t���CE���^��x�~+!U!H�8��^�uK�^�"�uU�}�{�!9~��g}���z�����"�,��է��78���$���T�����)�/7u9ҽ��
h)�g�)�˨��
���4 �H%z>���X��V��T�p������̭�|@���	C-���o��r'&�6-��o�҃���.`ʂ%�G�#E���fl�DZ��j*��zuO��aܛP���A����r��Gėj�6���-�yqZ�x���$����`M�+9&���hQ�4���z˛��7��Ԍ�6�~�X���X�;�Lձ
�W�j%�����+�����{�k�����P�: �v�4o�-Z�	ۇ%�_A'`v��O5��6��t���,oYknD���o�U��*e�C�4�_�?s�i��S��_�c=��#.<ǚ�[� N�ם�d�3�Ib�"��Aq�3U�κ����ҍ"67g��/;��鮊@�\	m4ht���^�_�f8�\��%���S^*S�`�	�|�0��u�%9�؅����X��i�M��_^�X��vD��h��^gL��/�j*q8��ym%l_���]`���+F����URJ��p\N�l `�a@X��@�2��)9tM��e;���c����� s`0M\��x��c���5�gN*IF����^�$����e��H�j=�3Zt��TQ>'��)QvI��7��#���0�nM�Z��~��#'�L�CO�8^O����ϼ5R��k�w_�0�~��Z��<9Yo
��H[B�G �G�3~��%�Pwq`�M�B��(ۛRb�K��c��f��[�b��Y����{�L�Oyd6qL]���G:E}�ڽ"]������d�����U}�o=���Vu���ۮ����2?m�
ʞ��	�$�]ʘ��|�p��P�iA�7��XJ`�w�H<��y)"���,Xl�$]�����}�el����g�,t���3k����_3���o��Q��}Y��ۏ�/�C��B��,y��l*�2=sCyL���nuS��{7h�jDGʐ�}��3{2�)'�Q����b������w�P���+>zg��OFu� Ē]6��~��v1��m�5][�FkA�����\�{J6���  �ف/uY>h��j�@��hNjǔ^��#��h�>&�7f�>�F	�̣k�$|&�e�}}�̓&��jxX�rbh����!��b���m�-�����
�"q��֍DU�)���$HA��M��26���T7~���fs�����_ҳ)��13t�h$i��ȯ���u"#�Fb5��(Qx*]OW;�c�9�A�w�k��	�WC�oJo��
�2�~	�lkȔç��3�Q�[���z^݉ �u�w�KF�c�����d]U��Kz+鴕��O?9"�ַqs�h�7�ְ�5�R���<�X�4z��S���?@Q6�`Y���텤���2w��S��:@�uǒ��w"�^5����S!)�<�ġ��=j^�~��0o+�>-6h��*(��\��;r�a@��vZ�o�w��}����a
������QR�]	���՗��cj�g�l:�?z�?�ԣ��-�_�mٿ��~�<T�0�	J��6���w�#�"���J�+�H�X�����Z_G�H��(��z�(y}>&-��	���J���Fa����N���b�,����m�c�ok�n��D�J�
��-߈��fT��.'�L�H��!j����`���%�e8�NA����5v4`��1�+j�CJ�z^�I�?$^\��0NE�)H��5���&���,��J��p]��?�	��j��,��XTohH~)@�)�z$dX`��	I'��	�s�	�!K�f��3����*��֫j�d��~X$��cҭ�W�h�?��k�A��^�`g}����pb���yt��>�o����0�񈣕W@R���Tc����>��(����}����֮
�<�v6J��K�ְ,���G��Dhy��"{d]��&���u�:��+��gI�0�;��oʾhw�&���s��ױ�����`�V���d�tY��%H�a�ɷ��5\Ұ��T�gVaZ�=p/�#�O%@���M-������G',�q[���	��6Yw�^b�����K�����#>���r�7�_z���0��(�`�tN�,�z�,�h�/���'Ǉ���U��9&G�[o�E������.'�<O-(2���r�ţ+��hS���¿����Ks��%GV��;+�@aglK/��&�r�����HX����{Vja<I�q��$5i�F�e��.����Ff�dNb����,�es�H��M=ߵ�`�2�h�� �ie��,�]��7SUA�8���]�O�ӽ�p�Q��G�XLC�lA�tFJ��1�xڥC-1fò>e��}���O)7���^��}��⬀����tN�<:~����Jd����j��ca�[r�1o�'Ɂ����������p(@�tHV�)�NAz�2诳��*)����#�
�8����6��5 H~i�9��&��L�R����Q+>c���F�/�X�$��F�
��tP^e���~h���M]�Y���&y�Ӯ<_��=��7���lD ̂B\�'� �Pa�CP�k-|3�(�BLvh.pxh�ۓol�p��m��[fUn�i�����nOo���"���;�@��cu�!���x�G.��]rE�v*�S���ek�I%樋@*,�`����:h/x!��U�XbZy�]��b��k�jyU5,1��	��F�Ѱ"��b���W�d��q0,nD_��^)���"��qb��9���l�ѹ���Iړ?ydێD��^h=� ���Y~��#�\R'{~��7£BGw5.L(N'
�ώ&_��S���Ɠ���U/\D'5g"�$�&�;�V�c$��������(�7�q���]�Zl�"�H�E7����G�7���5h��6,�5�ُ�VL\Z�4V,�{��3(��_p��ѣ�tap,�8
e�N�`�o��2|=��k�a\�O��Hr���{�y���nV�#���)KSF�9���	�%�T����]�,�� �G����Ы���c)�{���h����y�q{<�͂ؖ��U�T�1)Δ�֡A=:Ig��'�����0l<�<�����f�u6"�RL0����� -R>Pj�PR�"�̈�!��Tr����ĶR��y8!����(ő�'#�F��3
u9!�o�8<�m�F��؄y�L<_��V�8m�Ig)0����9u�&0�6*���fC\��i�8�N��uI!ۥEt���j7��3���̫�X�+� �N�R9��.���^�GI��h�L�SC���� �hv���(.*8���;��X�Z����wF'�$��,�P�!ݞĦ��G�Ā��<c�V��
މ�c��pPȞ��`�Y
a��	�:��h�Pkr�uVhV@����\%a�Y>_u���3R�D^��jy����J27���7#6��U�������&Y���"� C�:%������yj�O��)������5�q�;���b��zh�t��-G4�
��ݬ��o�J]����?J�C[�F7��3it��]-��!�09����@P5�g1��jq�s���0�u����z,v�D=Y��ꖎÞK�Owqp��̮
<㏡���Ke4Iʠ�l����`|��x��츌�ڌB�e�T�� ��=9�d��s�a��-Ͱ���}F�
6�*:��N�i5O�UW���R�J�$Ur-Fpt��$V�λ�Y�$���n�Wv���p�&��@�������
�ػb�+@F�Ҳ���v�!!���j@��À�G���
���UM�H��[��=_�+�-��}Ȫ���o����&�x��883.��?y��t�p,_��o�	��`��͈Fܸ݀�\߃V&�:�?ns�V���G�@u��q��d������{?qN�g��
kJsh�t�,*��Ҷ��:��v�2)��%���m1��0�'% (��U���HJ�)�zx�D�h�j= ��Tn/�A���WP���VY���A����� ��Gs_g�Xbr�^n�P�R|�n0���� y�.`{*��:�oSD;/f��u1<�E�!�f	��6/�����q���7P3M�6j�}촪�03)�Mw� sd����Pp�Cd���rz����J�� ƪ�e{�?������*�q�$<p!�Y#����O�fU"!kN�G��]����cFe��
a� F<�qvK�[U�pTe�j�'�o1��v�`�\�G,r _��A��N�_��I'��$�ML����r�XM5k!�&�fR̆@{B������+-}�%���-�?bM�k��)vV]�{�S�\\zyCЏa���1?�3+~�Fфw��{�*%��N��P�Opˁ�{�P�;�C����a������3�o�0�?��P�z=��*�r'��n:�o l�8#n��f��TIdyZ��@�2�Y�O��l�H�}uG[H�؃�`^����I*�F3c�j���v�f/���?x�%�
�ƣ�nT�:�.W&v�q3$��a�Ὅ؁ ��6� M>l�4���Ep�L����ʥm�d����}����o]d�����(D�|9Nd9bY�t3�{�mPZ�.��VP vw����ivj�&�le��B!�.��v�����+8���.����9���fXlxVHYEB    2889     400��X0�q
	�b�3�Ǆ2��d���]��� Y�n�n�'�r1���F΄9`}
7�k���!���$�<��� ���[-�&p�2����4�4��T��&�,$�G���lZ#D_����Ö��05�#*��G3���Z,�����B���4�ֱ��#�o�tM~}�YB��g�[����X8R�R�x����^�WHm��y8T+��),��k��[,p��{���@���_����=A�`LM�����4�X�I!3I�{_�s}p��{x�דx)jD*BB7"���u���V�ڐ����	n��[@]R�������H�V����}�)��ϲ�;������\�f�C����K�����Qv��N�P3�*�3*���խ��(I.ޅB����<O4�_�ܼ��%/���"�$\�3�ۘ�jAU��w�ǥ,�k����Д&-�:5_���vO�`,�b�3re!���}��9��29j�$�\�ec3 �4@���qX��ar�;gBψ�_�I�l��q�_%��I�+�<�ܰ��Q��r��[��>Jk�_�Ҏ譀|e9���C�D���g��b�[g'�&���HO�|Y��Ue wx+�A(WD^��f�b�@!'ì�iW�6�򨈴e��`��"�Kv��cl����|��D��R	���2�D4{��|Q���>~"���%������9�
��[��Bݛ�iS�u*%D��8��E�^�eeU�(���c@u���ܓf��J!vƯ}�j�Ӛ4Y(��+!��F�uX�6�1Sip��F��k;��1~l��`��h)E�]�Dg�4	gW9V:�Q���2K�h�kԯWՍ05�KB�8���7�D�2��?`��O�j쇀�,�Pr��B���|�����W.�^
z�7̬Cb�J�EYq�Q��H�]b���ϝ[�H���6�
���x��B$>v�V�:�rw��s��Œ�������_���gW��3ۆ��7�Y5�x��������wD���/�i