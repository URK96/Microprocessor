XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���&�V;�0��8'�W���y�Y�UQ�[�?q�s�/�N��I�v�r`[i�� ;�:� �{����71�4``��V�����d������g[\�7��R�HwN΍$�:Db�c� 0Y�Ж�~5_"/&���p�H� o���b�FM> �� �q��JmT\�>g��]��rޯ�����`��#��8�q��� y��03�t�Ȉ.�|ˊ̪��L44:�C���3�;�H�2#���%'int+��p�t��yS�Ά���בMe��l�0Fx���3o �S� �9�5rW��}v��~O�9tc�<���f���|�Bd;$����?S�~wl��` vr��r2`u�����Y�?�����D��)�(��L�:sb�Ok����F��g9�9�����S�d��%���_O�l�.�zd���amf��C���ʅ�m��lb���g��G|�n�$���6�KZk��Mk97Psǭ�K�4c0o0���"�m	gH�7�^��6a@/[����.G�:����0�����S���b�������۪�,��-�vfaG}	�y^�����Ԧ@�t����H�x�2<��6}
\H~J��:v5~4ɡ[��U	�(#�M���f�=�OKl^�9�����O*�\G�tL��᪪�wz'����j�2Xa�?h��\L2�u�@Q�l�&��;���Y��_J�I�=��1�+���Qt�*mpd����z=��ʦ�������E�Ez�Oפ����n�%XlxVHYEB    3c92     900��2�i� K������ՏZ�dd6��>�,n���ZVcy��q�a�RAϕ�ޑ*|�Y���m#�o��.r�Z1���p2����Y�%���3���Qr����r�y�@���d��2QDUO���b���{�xxH�D�����Q�vY:���@��f�i�B4�O\FF�u�m����� �Ck�S�����6�pG|,=�5�����p�}G�1h>&U~��,���f����W�)3��˕�=�d�'�ߐ�$�Å�zk�N��с#7��F)�de;�0iRƇ��y3�Ƀ����~m����~��0���ɌȠl���q5���z)�6�y7�A�Q�y�;��m�fk3[���ڡªK�ҫ�����DC�f�{�U=`��1�v#�FE*f�!c���G���P�!m�t��ԋ�T��z��]�iq]�s�^�8	������G�����yΥAg�1�����`�FJ�'���{���y1�Bg�/���pT4�Z�5/�S@5�q#�}�	۔vc�L~���U�<)ˡ(g�e�m��Ax��$�r �.@�,c��¤��C@�̦�Ca �]�z-1Y(�s0��� }w-eS:�k�D�U��n+���}���!�yGY��o}��p
G�f���3����Egwt�=>���a퀤��'=���1e0>Zq����qR��2�!K��D��MP��p������#�M�h7�zC,L�,INhL�v"|p��ég�4�c"{�L�i��1\����<^S&'�Ή��[��z�B��WԲ�0^�8S�bVc�T��>�e��I�B]���I��'�s2�=x?���9W���"᷉�����#�܋�7����P��Lvr_�, �MN9��{��5��m_�����IkP��N���5�J�t"3'-�v�.y�k���` @�Ec�����Lw����zYA��逹l���T�7�x�@�]M��b��'+弶��K�&&$b'S#6���G2��%�~�ci�,���b����q`����,�Ә�����я7`8�1vߌ�5$� ���^�c��Sb�0���7F�Ƃh�X�g���Ly�k��
�9���qHj���0����Xb]nv��[p*N����Lܜe'�Ưe�P�؊N�˯5&H4uC>�����M�z���` ���`��g"e�������w>��O�K��`���̵n�
+��ZI�����f�	�pѕs!�Pc��v��Iǲ�nI��f���Ҋ��X���K��w�3]�y�B�@v^Yĳߎ�,RY{�#���(�@����R'���F+�Mv%�����Ը�?�z�<�qHb]Z;V�%��@���T�nGC�p�Á!}��ԡ 9�r�]Y��'��A?��e��m8S��F�x�A��˙���xf����$]��#\�-S ��DT��q��R�V���$���'ԛv�=�t�e�)��X�C�jU
U�d�Ԁ����fMSa�/;>��4��*�u������Y�-s-�O�q�m���x`ߴc���r!�յ��F}j\&�4G�*G�=L�%�׋�����6�1����]m���qH�<����왇p�fu`�?}y��,�Y�u����Z �x���B��s�sr�P�HB��yBo�?���ITƠ2��>��T���<�>H-��q�:M�R�v��!�Ħ
�2�|��h�(OM�iچ�_�$,�Y/o�Vd�����'�ky@"����qY���M�E�aj�ǘ� �ϙ��i�D�l}��	����uKפ;p�g��[�j����u��e���=��'��pu@Uf�L^���YbȄ�m6�UOB��"��E�����}�tŞ�����`���Éx�Yw����YoXz]N��zRu�U��\|���1����-l������1Mid�=�o��g�c�P�p҃����z� �`�Y�Q�-��\��]J��s�;@��W�<���1S)���`����г��	OW�f\<�3h&��0v�����-\7�T��9N�mg/`����<-�@�m �6GcbG-�C����/NyͻV��فjI�V�7��luq;�J��nG����%7��	��7�_*���<����
�!�ok3]���1	�I`��x}����}�D��Zi|�5���!�����N��^,,-��˷'�Q�G~D<$�p/��ݫ�pVr9������E��!�r�U��8�qۄs�"��-�0��.]	=v��<1�eW��I��IR