XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[�%���Aքʾ�,�繸��� (�I�@)����퉋���o�77�ܚ�ݧi�Ur�����9�0�ꆪrbt_v\ �/���=�т]���N�1��|��=���u� E�LwJB�C�Ȗ��I �q���ic��EE�ޠ��2s]�  }�Ų������j�y�W1D��5k�Eiv��Ύ�`�� �4�BQ1 ߂K��/*��>�l�UP��$������h�x���N	�%k���yR�&��[�o[/ߟ���b�lh���<@ s�2���;"5!�2?�%�={~�`J�ÕȂ'��㠲Q�T�)��t�|i0���e�T���/�#�0`�s����g|xz���k2��
�v�����!7rf_���E�L�C�x۸�c.�S��]��#���_g0�]��2k�8B0��T.�c���Kb�1T]Mt阁�3���%�50�CP`�y@�l�������;rW��-ǗԵ���Y��i��H�����g�o0��?�A�Ɓ~C$�/�a�8�9�_��#�������N�W���.����Nd�y��@��<%߯�";�.rx��G�������&p=`�;	K�7+R#�S���N7��Ԁ�J׭�.�7�5��UB����F;R��W�Y1f�c�񷷕?Vx<E*o$5Ԫ���X|��B}���V1�% �>�r �-�`g)0�OW���:%����{Dq:- ����m�L���>�n�H�i�#��@z� �Cָ��Y_�(���XlxVHYEB    2863     8d0/�Lc�s��76T���(  P!H|����!P�+&`�ը�<�����`��H���!�)���
�p�U���u+ͮM�?0wyE�K� ��������%�,#x
�Uư}�ʵ���aL�(���f���˹�So	�E�wF{���s���MN�U�b�8_��~e q<.��hs�"����ä�K÷?��#��moH%�����ַ�Q��E�}��64���@�F���uùB�t�3s��{������@��{��ۃ
�'��Qꯒn:Zɴ3�`s7f����f�V/�#��D`�$Pkv��x Z�8U���j�P�<7C��k�
C���~�LΌF/�L��W���M�I�۠�n���s=ȺN�5U�J�N���@�4�l�9
��2��]�~7ħ����Ǌ�\m�Cjђ��w)�=���둛N����Kc��4U���O���0����e��v���8	0���ʁ�C��l��1���O��x�7mǛaW������]j��N~��_~F�f���s=E�q�p�Z�5k	���Ŭ�J��s1i��?tE�R�-��m|���p,Y�T��2��I8�	���H��~+�H����sZ�&m��ē�*���Ģ�y�����9F;���˯6��-�`� "�� �
���D���bd8� �GT8�hr�{���;2-А.���֘nt6`w��pB�����R�����T�heک�*�3�!�����6���N�W�Զڃ�M���Z��}$���1��9يz� �� +A9>�>Ｑ�a+�����f:"($��SiI����s��'����	��e@lw�t���wR ��S�X�`��'�*d��$���A�xɎ��*�Z[�*)҃C�C�9jrc3A4�G! (Ifm�Tk��;�ws7fat�.�!��&��<��m�R���T�$7�?U��P�U��g�w1�o� �?ہT��'��
b��uPy�;~o�k#�H�=�R]%+�]�{�G�BwK���$⡻��rS�p*NΠ}���vu�]�9.Ifog�3�	A3+r�:�D�G�g��Z���6�fP�_i�no}��"�@�NI�G��~);��wG�P���euT���7r�l%�+u�b1�9�"4��g^��a�s�{�g���
�-
�Dc�$����Q�T��W�����$�4����p���7�;��ϼ���ܵ?�8�׏P@a{�]x$h��#�mcChvՈ|�Ͱ@m��`}D���<ܱ�ҠaUT�I2g ��G+��!j��ڏB�3=�_lʫ�%O�N����K����,�[��\ k &���1js��t�k�d��^V���,�}�����L8N�#s>�L��� /#�x��kW��u�^��O�R��@���ڴ|KAP/S.�+�0��LtF=Z��1r6��$�Xᤍ��.��ϕ@����Qn,���\#S��Y����Dc�H1�!U!��.��LF6�
`�{��b�J׆�4����^�����5�z�3�m�C��l�DD[ ���!�=����(婈����F�+�_kW�D~7�դ�+��Q��^��;"y���+���-�:Gи�S\��&���B�I��mb[��h�ގ�ڇ���Y�J	<HoM�o�MR�;�S�����&��=s߶.ܒ|,��	��kv>�L�r�NK���|��;�a]0������e�����i����aB5�n����;k��B��c��R"]��ٗI�/�)�����vk%��A�sG�ߦYɩe/	Vp�f�j֗`k"���ܢaZ�1�"su�=ۡ���z%����Yz	ey[�d���5Y�e����3)�#�b�(E��$n�.����'#:?��+���x��� 3(AL���xG!H՟,��!�e��dV�H9n.�F�44<�^�꽟y���"6�a��(��gqA�س;4��.[�9k�D���R��Y�ݽܳF}������P1� �U�k��3(��)Vo��,|[������?Қ5N�l�h`8[�᳕��t[��D��~w�$�#�`ŀ�@Mz�F�[����oV!�'<%����o�k�>,�O�.»�c4���8�1pg'|���KŒ7�K���=UdP	q�Q��Z@gm�:��M�?�m��r(»xa$�O辀e�c/��7׆ѓ�]��݈�\_�)����T�.��%���B.(x=FK��X4|a���4�$#�݃�����r,��vO�R�