XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���V�h�����P���¯ت�=��)�w:��{��c7�*Ϧ��X��r�������'�d�%�V�Lc����Q�K&u��l���a�<+i�7y��8�r�ނ�W�&�2�kMs*'�}�܃��d�"OP������+QP��(oz������=c��f~��׫���{uW�t�di�԰D�,��2_<�s��a6B+�q+�w�-��Pܧ��u�G�z�j�ORU��u�B��|��iLH1!-{�/�ip�ÚǱ��>iI��h���b?�I�Я�����S&�6����Ř'�v��K*~�� ���Bx�қ�8��&�_.�e�Ev�m��R4h0D���j�����(��]D��b�I	�|��&+��69x��H^ �G��iUԞ�aK'�]��"���+�Wj\*���M&�H	aDo�S%_�_Z��ʍڰ(�^f�{#����ХZ-�頠����j��nyi�eiȬ�ms����Y���b�LD* Q�ݚ~�RFp*x�Vi���/�Q��zT�|�K�_�ĉ�Fs:n�e�g��y����Qj�����(a���@S^�;bɜ�F(�O����F<F�"F�l]��NƫSx��}��Ăo�����o�?',d;�a��^x��Tt��?�\ћ���
o	�a�ܵh5a��lY��,�yl=�裖��)-��1#Le�@w�lQXEY���de��`�`����u�q4x�\��� ��q�w)�65���>�x���t��K�_)Qk	XlxVHYEB    156c     590�'��Qj���N����^8�,YͰY���MP|�\D���Y0;3�v9�t��B��1\�kϡ�|+r�ԧ4���7�5:u���0�y�Έ�G_ɾ� �K����Pp�;O�)���i�Q�>����������4<���?��'4�7? @��6�C�(�Z��!c]��4sw৚�'ȸ+�D�'��@��/傎�l�z���,Cz4s
ȥ���B������PCW�5��+E"5�|�����&[Nk>��G1+<I���-�&����"��'�+����s|�=4bo�Z�&�B�&Pw1*Ct0�1�1R�x2��T��jl�zg���iW������/y�,��@S/#�9��s��;ɒ�+̮\��L�,\�4�׻�
�0��ms���$i}�2:h�q��X{�2[ؘ��u��{�zv����X�P$m��,�VIG|"��JP�J�G4�X���;����T����A[uh�Jf�7)��V��KΔ,�E��Ag�hZ�,��LF����;��-�(x� >P~ߖ�5���8~!������,��@��d^lW�	}�v��U4;�o�B��e�����#q�%���f;bi#��E'�w3����J��n7tⲧ��\����AMq~�I/-���c<v���r/֛{	��[��X�A�PK�ɜj�� �C��H�7!J�FXo��+��˲!3���krb�\u��=(�*h6qG��<e�fұX��
-��3=���u%O�`���D�D���ޙ�g��_�ҵ�]����Vf�gf��ihŇb������u��5�O
��h뵽]W���1'��Z�To[��T)�������%c���P(*x9E}����O�ٖ��W�}�	4�&4WԞ�ʔ��yI���0ɪ(�B��E�~�O�j�&n�n�_8ֱB�#O��>��#_�;E}��6���<JS�+s��k
��}<�׷Dw����{k���4�X�@r�*�*'��:�	�V��.�IǦ�C�=��[� W�I�k�R̞m���h5�`D$n,�U������)�Ͱ#}�-7@���v����Z�� ��Ʀ9�>[�u{�\�m�W�
�w�]0A�fl��p��̖cp�\m_�:�B,�Yiz��".�:�8p]���ex!�+q�U��'�J�J�\DHr��6]^��y�r�E΃��4��g��.?��,��"���D�	��ʹ`4,E��\~4)���O,C	�+?�D�7)��ű>��A����5����]r�\34f���«�04n���0/�0'X���� ?bԟ�h��v�|�� �ě3-Kpr7?��Tñ�XIs�?����us��H������x<ι���e��\!��Q�TGd[��.b��C�