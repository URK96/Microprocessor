XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��޵�+��Q���y�K�&
���Iz7i�C N�s�rh*��%`���ݎ+��,f\������_C�*�=}�ņ��+�S�vM��Z�FXɘ�$�u�!�F�Ӓ罻"����2��}+o�b��r���rx�hi�@�j�|�v<3���G����Ga�0d�v;7RN�A֚��U�*���n�����dhK#�u�p�|���	�N��5*
����Q�������U�e����'V�SP�*�����q�q+�C�۰�H�0ju�!�T�A�na*D I�f��r�����M�%9���|���Xi�3Z�Y���3Kz�Ͽ�?�t>Q���&B������e(��a�(-V ���"wf�
�
��%�_U��ܓ������]�j�O��$!
a�����,���B�����y���tݱ��-5I(�0�`�0n��2���/a�l�/�����ٌD:��k�Ck0=I�e�� �봴��\2G5����lN�%�}��0��2Kd����P��"�*º7���^�w�a�?^ĢB�8e��������$r ��d�R[������9�����{JÔ��!��(!+z>�j���E��/QG���O��z��S��� p����E_��[��׶�^.�1�s�E��"�e!T6Wc���&��{�j�Ԡ|H�n�"��F��M����<n���E��2R0��Đ"�&޻p2N����kׁ��si��HG��Dc5a305kf �� YiEx\���{��f_�0m*����XlxVHYEB    3c92     900�.���zd0Mi8�^�2[����XS,E�GWL)��P˦��|�L���^�����kj
T�2��0|�_�|ù#:B��&P�jq)���?�%��Y��3@@&V�w�UsΉ�����V$��Mo)O���?����O0;�n
��R�`�o5�v�4fs*t]b{!�i.��(�3dJ ��z��)8B�7����n��{�H�?�m��kH�pv���Ϧ�㠬��YKc�a����E9r�vdػ�����x�z�������+[������Ŗj���~N���)�(�������	�Ϥ��^J5YѨ&`כ�l�}4PqI��`�N��sa�ª�q�%4��I��l���>l�h�r\���n0�ѻ��M��Kcܽ��$ʪ�=���u�o0Ǵ,���o���F�&��
�5�*��v0�>]�zc)�Է������Oa�/bځ���,@u���j��)������1���u2��M/����;�VM��hn�	{	�����o�m�b�:TpԹn+C�Iv��ǌ�@�[!��a7M�B�#�M�J�����L�vC_��噗��[k����N2�X�L�0��wX1�c���+W>I9vQ�j�ToWor�{�B.a��y;�v'���i�w���+�2y�V{<c����	��B��k�i�R�č�8�3�/�=����8�4۬�x�s�ؔDc�qp�;�02�#-Չx`n���~�V�F�R�j6������=?�m3�ә�����P	"�/�T��x|�O�$��/�y��
IUe�L�vQ���i�=j:�^�^8�]�Dⷞ��`Rq�����[�)V	�+J'�����C�S����sq�y�HE
Þ�X�ߪ=�{*W�q�K��"��Pt��z���pҩ(l;�ߡn��9��w}s�&�C���E����EV���8�C(H�h����Y�t�����,�6R���U�"m�6kjM<�e�U$�5��֣���E��?�������}��\c��+t���E��oV%�LE�ȼ5>Ƞw�3R]!���Ġ��4=�Y�!�w�q�4�������̳W#�<��0���qH
�Քɟ�ڮ.��_���X�=ޢW-R�b�@�T��F�$:����ūm&�+�K��tY����\|�Ub"������4�Zy��������xl����M�ye�ќ>4�*� ��<\�.X���~8���?t��}�`zdR�� G�i��e�� �N��t���2"���5%��,w"Z��`�g���V��V_�����_��v�t&�:�-c}�O���eP@����������ex��$��A$�x)�i�O��$ygMLF�ʮ,�߃^�X��,�v�<7|��/����"Y}9\�>/�*�m�ξo�i�ʁ�#�Q��J�3$Q�k>���Й,g��\
q���ڴA�_Ea}�00�����t� \�<������B�s���i��@����H���½>s��y���`�1̎�(*����!�� �B�U&�ѧ�k�ػ��{��yj��pI��z��ܼt��0�i��Ӷ[�-��a,Tڸ��P��6�fE�y_L&��<�����J3hX�!�Cqw�n"͞���yIB��o%�������n����6.�'�i-�b���t��ے�8�[3�5���T�/��`���-Ϻ�N���)��CF�?WU�ȋ�lt'7�9�?S���Т��P�bKi�����O��׊%F���Ҧ���4�tN4[]jT���7/��<v�	M ;O�/5=��ܧpEVڋR�_@ΐ0S��L�C��ї=S�/:���	����eƍUF<p��$��b�II���XI��v?�U��f%`��Mft`6C[ib���Q�L�<�$����.!�K�Ûs�zH���M�am0���c������	�8��]{p�Ik��>Ge����3WAM��7ߨrs�b.W.����C��Ĕ���?�b���2G���u��R����'��`V�QrF�(�N�:d�~��Y\��IfC�`�����YҀ��7�ƅg�*�n�ac�3��䥢;6>_����ʫ�������~;��k�����x�f7�~��
�sl��k]�2V�Oq	Vew��'MW���ڹ��`�J�����#�|�k���Uw����`{��"���YA��(��u�"�����&�)�-�іgM�)���q�No�C����A����h����Og����	����z&�Y��ܿDh�eI[�(�fګ>s�`�w,���z��|QrG��Y��V;