XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���M�6��}���ղ�2����R��w�d�j`���eD�B1���VTz��ǏS92R�ǳ��[�"��mk�F��brU>Bj%�&��n��{�j��މ`qR��K���Ѭ�FK��y�$9��>�vD	Or^�+�S
�x��#j��qz*��J��O�B�S3�����$��7��iІ��#���M"��xH��ͤ��R���zm�z����E�, p�
U�CW�1����9 �[8�ה��Y��ri�׉&��$v��+	^t)T���k=gv%�btW�J��הY7o~ ���p*��W�&&��V�Y�-O*�H&�GzM���QX��غ��x�Y�;$�p���W�'$ӝ���J�T�L�	������U��s�y)�A�5|h.�)�)����Z���Ǉ'����s3��� 1~��'�`���k,�A0�D�'��a'��y�s譁�5�U����K�C�uwi���Zf�;�o��De���G���\oֻ}�������=�����$�E/&N��˧A�њ�F)1�q����Q���Akh�%*
1�z�M�$�%ڈ0%a쎇mN�L�{�4c�>y{�$�ٸ�A�%D7��
�+�i�v���1nӿ����A�Yl�-f@�,P�荩"�-�%0��N?K�i"�%�| �&��<e{�GĒ�M��` � �=���"��Qߒ��:kƋ��.��_�xoh�n��3�A�����/���r��hE<�PRg�:>L���,�Ƞ(�
��]�e2���;z�XlxVHYEB     b8b     3b0߫?���&�Y4�ޟ���M�27T1�Z7��^�R����Ŗ<�.ֳ��!�����n��eD�r�̰H���W[k��]� -_�:��o����N�����/����Ѣ����ރx�^���ս�+���X�FP"���VUn�tu$���vmm؉���V�K���Z֟j�e	+��jYȜ�}�ֳ
T�?/�(_#,u��r�}��e���)�}NNV�0��]Ғ�q�{�CM�kg� ��j�q�H��Q�ʖg/a-��c��s���u���@~#�ȫ�B��.d��k�A��|[���3Җ�t �9c%�/H�݇�wp��z7��c�`�c�����e�u�����M0�O�0<&V9�:���W��*�qc�����3�� l�(��<I�)���v���8GY��H݂禃{�f�
^*�I(�����~�3zݡ�"�n��m���Ʒ�I�)�NU>iA�,,5v��A��?�\�B|�H���-/
�Vɝ�q|��I�e���v�A�80[�S�ptĻ �D-_�_��o���꓄nN�+nҮq��2���cۍ��3>�2$/w6��y)�N��4�!䆖�����ez��}��Bs�V�O�X��7xr܄U����lF9�Y��cZ�X��+�Q��g�`1>Zn$Mz��&�޵3R�U���(�{�X5S�sH�+�V����Jz���������Y˻��i��t;��ϫ8d�3�tPT�Q���')d�p"�e`,�1�6�f�ׁmD��ɐV��Fn��bh�8��D_�eb(�C���B*\��'��9!�Қ�%�뒣�lдk�c_� 1������7��r�A_#�����G���I�iJ��2�C[2	ֽ��'4��Rs�a�JL7�Dx�K~����י�i�:Q�b+Y����C���J^�V����f�