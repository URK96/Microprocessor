XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Q�����ݣv�'�X�����"����O��G獘J�g@E�����_-̻'��t�Q���TS��~�.1��m4�0!2�۱����ۉ����Mj!�X(���������R����6�� ��uح���Ɂ0�B;�F`���� +��UvN�zU���7���x�]��iڲ,7���V?
�9d��9=�V)�W�|U�i���oiR��>Q�8I�����hH�l���������n `�W�+�z�! ��+V(U���s��FS.�X�-eV%�����&�^�3��{�IQ���c��n*k<���S��6ƭA��	�"��2c��͈a��L4���#��0w�WO��d����:�x���� ̿�E�7g�롵�bۜ�Y$V�<PO���2��G�N� ���	.�O����ϖ��t��M<�ٱ�r,�{B��g�����yf��t�MĐ�	�cP��.K1�;A��xX�+U���j.�B���� AI��?������g��5,��I.�c�>m�ue��	�]5�<nv�1]��r�'�!�XN_~��<K`���2��N���u{��	�`y�"t���R���19{�����;��ce��^���㖡1C��*p�)M�14�j��5(Z�f��2I 4�C�Q�#�)����8mŋ���G�V��щ�?��?H�嚜@x�s7����\6����E�-�d��u�E�)��4@�<;�h�+l��ai�f;�	�ŴH4��+�u�|����XlxVHYEB    3a1b     d40�}�~�1�ǻU��bD앧��9��5FE�3���ʥr����"R�Rkc�c�S�=tG�`������Ϝ�y�۰u���u�Կ�dHF�G�����(]̜��\�DZD�K�Ie�c��Y}ͮ��
�������Co�it]l=���|�r5���8h{�q���%�%s!L�!��_�\���� � 6��w���/�Ż8y�6��j�}օ��7��mkUuS������V�������IM����x��q[�����fJ7N�=6�[N�ƥD��=o�M�����վ-�HwY<a�8�5��1�x�\oA�6�L� J�-W� ���O��~C���*S�P�]��Mg�ϢDr�[Y�V7��+fŏ�t����H�Fm��m�^���e��P����o�E.Cj���~
+�P&	�G` ~�. i��?$�{�ǌ���2	]��2#�EX�i��	�&����x��c|��	�)=���J�!�M��ǧ��-�-��Y,	k��%��->6C�=&���%7W����U� ��t�P���J8�]fQ`Uᰛy6N�{�v���ս��7��eLQl�Y!�[�1���u�m?[�W�2�O0ţ)K�A�2=a�f`��1=����jWL~.`�W]�8�f����+`j�f'ł�H��O��BlI�2��iB��)�p�XmG$,�\6h�M`1Aj��;���gNsbUz�/� 2c$��J�^y��w�
L�1c�ha�P6���{���go��w`��b�`�]Y����!�:�r��
�p(6�D��;a^1�ݑ�ц�I�"�'o��&;#�¦����*$a�R�oG���J�w#�ɪ,�?�t|E��<�7u`����3';�C��x�q�� ��pY���ų{6 9o�.�*z���" E����#..-/��h�D���6�sKC\�T2�4]+��`���Ì�ml�P��:{;���;rB�ń7��ۣ���)#��E����Z��p�[a0�����aZ��gϤ�wKC���˨aM�è��BL߮��Hvu@�oe�*�/������1죸��?��͊��"I%�_h��Y0���)��D�v8����n�\j�_(�!�8ow�/���,�����',���Ҳ�აË�e��A?���׮:N5f���=���t���t�����wj������U��` ��o����*��Q<"�S�$�4�XO>��l��D��@��`�P-��Ii�ɨ�S,
�*���ލ�m��|Y!�f��!��a�d�
���4ʰ��7,�p� ��#8�ƨ��K_L��`Q�Sd�K%j�G��B
�Y����-��1bؒ6"������h�}u��U�W�kئ�3v0���Q�!!eE-�Y�͆~�d�'��V��l�)��I�n�Da|���e�S�S�Y;�m<��+��<
�-��Bы���¢��ߥ�R����h�`�������l���RרV� :��E��]�Gg�[��2v]�� 5�*�Ŭ�-��`�3�&]���1�S{����l�Qo�D8l}y^�Ql����7���O�e��<nkh�5�S�q/�k�2$Z#U���&b�0��62xC$S�ǙH��(g��0���vT���i`�����B�Y��`Z	�{ĝ����� T��ֽ�y��VL~��>Էy?������K���Z��[>����6�2!
~j�1_��]�j�",�X�R0���I�������1�*�C��$Ѫ�k��Fg"����9��J�"���o&gR��y]����f͍ͨ���X/�Q!�^n��P�l	���F&���CZ�]�Q����^�X�.H��I\k�L��� F�hXj��Z��h�4,�BkC�?ZݦVӸK�%2��sǆ��i��0"�~����ͯѪG%�����!����$��-�׽��%�Q잘n
���'�ˊoF[�L(0F�����?�$�4N8�x+)�,�������\�V	���y�nY��4�=�VD'�XS�+Tk�!8_嵨�����Ά,���<��SJ �����_�|��,R�rGC���׊���Q��Q�kʖ��p{�Gp<��YUG�zB��Q7� �/���^X4����x%�d�t[��p�w�tQGA��2�4�- �(0���4*����sK"c���9��	�~��1�9 �N�#ǉX��LGfﲪ�i�Շ��U<jw���Nm>be��������*��A�f���(O�8L�*|� <L%��iu��~���V�gKeW>�B���N��`g�NFXC[��x�r1���EL��_���NK�b�C���9�n��e?ݺ4$�ǰzq�s~F�ťk"��a�%7)�_���o�[���m�u�wf�{k��N~����	�c����=(���i�[D`�S̬��O��w��1�go4eH1q�����|�)̕<!��oh�W�[ѩ���Rv�eQԇ9�o�l��
&�h�F�4�R
����v<.3W�T�<*l�ی�L�Қ�%�PlTj���ƙJ<�~��-��-t��vN�"4���ǨV���U��y�ƨջ�� �׾�{����Nl�'r����7�	Ӭd����d��5a�W��4cκ��.Np����R$��
]��.�l�ͺ�~�~�=��ܪ|�����|(�q�6�I_���:���q|e��+.d��)g�W�Mƾw��h'N�qIk�W���ua�cGx||��\��0�+~��S��eH`CI�]�K&���D�0�\��$�J���p�϶7Kn� �[o���H�����'O����/)�@��#hut.3G,�6�n��
3t�r�wS�,��"�}lv��M�-Z�a�iG�;����g"�p�P�~Wp�|���;����V)�H��s8��x@%�ݻG�8��Yjj�n��]��L�	��bx;W�Ѭ�P(c�G�,_`�Y���j`��:��"H�a���#��>}�@M�����5�ve�:3F���� ۵уZ\���\��I~��~��D<K���(q ��D�m܂Q�����Mmȹ�D̦4�ֲ���o���3av�mٱ|��I��i-3�gC�Jd�S��[Ch�B����mppꂱ���羲�ٍ-�UV��.���6�yxZ�>q�x	�Uh?J�[�Ǜ�K��N7�O�X�B�JC/�F��\�����F����#�w�k'JV=S�hȆ���}��9�����8@��,)�����`��+v��\�9'$V��5S��s�8۱ݙ[��H�8�y砬������X���L�jR~~�|��U�s!�ۓ��"�A][�>��u��A��=۴��Ӗz��Z