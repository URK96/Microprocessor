XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����u78\9煮<�@r2#s�Q�ҋ�����6\]F�ME�]��b��;��(�o���]>�U:���
Dh���:Ë�d��*yvHh�_����
��\��+��
�S�Y��d��0��W���#�w]x�#�;����jG����ay x1�8W]��4Xp�.��w����[��e�?���ӓ�����v��wj�b���)�@?vO_z��$��	�/���^[ֵ4R?��U��PQF�5��k�5rxVQ��y�61�@,%Wt0<P��#��ڠ�g���ϛ��<[�[�Z�O�뗶�jV5n$�KN9-I�E�,k�_!!bDrF����[�;Vs�݃�����^���$'�ji F8��U�-a8��9�fO�z9����_�9�;���mj0��rp���2FO�qV.tF�@GwSK�lM�'(s�	�ĳƓg��n�hM0ZG���4g�R��:���u_'��;���l��tQxv8�s�V����(��'�m�P�_���v �#����7��S�%��Uπ0d�wk��
=#�i7�WZ`D8����D�.;�V��/�.�(lt��YE8�M[��J�Q�OT
��RW%���
�N��q߹&
i���Giل�nh��/��J�8�{�áVA�����^"]�ݓ�2�-������=N'<a��Fz��T��G���f���u�?�v�9!I�E�����ىv��9uB�����g^.K�x9�6�+����S�z/6Pb�.�k���J�宜g����<#R��]�f�XlxVHYEB     686     2f0�!�9g��}�+Ui��{��6����`$��pp7S����c���&EȞu������;�V h�M�K�֓R��<�\O��^ˏ��U��_U�/���h��rC�@��Үy7W��^�*_��5R���~v�Ln����|{=�;�v�4�-����[`�U�:"�=�N)J�n�rg���ã��0��iK����� 5�7�Wm��!YG�����mU��B:o�@���4�I_W�q�7/@�����
�K���%�P�%�+_JΤ%zC8�Wt�4$� y<�4��/���Jyb��'��{z	��]i�AA4B�4�Sz^�
� ��������TF�u!�}��,��pHy��4�5�
ɲ���N�L������yߘ��P��Kδ��
���X�V����Vp.a�ozw�-#��5��$k�y5kK��� "������yfI��Y��}�3�w>j�+����	�8�1b��#����ʢ< OAU���0o&��X��>R)��n�8$u��蠽)�ںfu��:"Hn@w����yYw��P{�8m���� �BDN��t���ȵ׮�{sqaq7���8�.}y�����@1��o�����Q$�_ �|K5�*y��ej�v
.�ԓx����'2؃K(m^ �p�x�"a6IzP����ȑ#�rGYc����1 ��([x����|���k��1�`�=<Z�r�:"/�V��cAt@���q:��@�hkN�1�Ĝ,��z�C�~~I��.���7�