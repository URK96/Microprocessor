XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3ё�l*�GŃP3��{��ۛ}�j:>�� ��"�Ӟ��oؿҗ;�_�R�Eg#Ý�Pˆ�ǝ���܋�R�HWWX��l<@�C�zO6�e��57��q&�'��>�������
+�|Y���I���/�t�5;����Le	nd6T�44�?I,����m��z�A����?�'�-��PG���})������?���r�Bk����Ω)�c��wo�4gKhaxZwV��Ч�oްeb�Z� �B�����=�|>��AA�|�o�_>�ͽZZ�>CXLeQ) ���l-�����,[��i�����!��,XN�[Ld�uSW*[�h������
�ۋ�I\^�3�����]y��Wĕ	�]�'�˔�it���#�3�3�+�H��s��u�
�k�+V7����������f����w<�G%�|�sn����OH�jG!�P��(P�I|7�P�ZL�n�,���!,�TQݤ��0��;�)�kF���H���`{\���N��W�)4]O-֍M��m��X�	#�	NX�~�H��^��rWL7�y[�!��}V@ʏ3T��Y���sX�T��}�JВ����&��oM/�e��Z
��OL'��s���	.�D��"�P�.�a:�(Q� #(/r9Y�4ׇ���e�BzB�K3��0�>��(���\`����������Rp)rZX��^����%����j̙0��]p����H@��*��ǜ��	��L��"K9���l��+?R�Sҡ%�m��DB�F��� �XlxVHYEB    1d06     5c0�y���M�4���H��?�(B�^F繤��BXd�ݧ��>E-+�O������Ґ���i�Q��1옗��.HB��Zӌ��o����� �	4�;�8Ԃ��׭l��0���������3$�X�VR47�N�lVo?���zXBM���k%=��2"Lӷ��R}BFN��*���	��5U����oE�����6�o)L�՚F(�J�,��+��с��Q�<_�X	��
��J�F��nH������Aհ�̼�Z1���D(X\hs@����;ڴ��d5�#�J��:��+���m�3Y�s?��Qd$*u�|�ۻ�^�Z%h�U�����=[�_dU�b�=���{�;^�w�֜��r��8�Tw�=���3{oFI4��9$7��u\6�M�Y	g�r��36ݛ��[G��#o0������$v���{p����1l4o��ӝ�'>��Ċ�i:(�U�*���� h�AG(ܜh���|59�t����A1ټFW��TA�Xj�f�a��Vܥ�;X�w�l�9T&���]�R����D���AM�u��r(��F���ߪ�����T��(i@D��%#����Qן��m��p���,��pj��>��} ����N�@�8JfQ����!(�&����oQ���e��o�����c9�������T2Z��¬��&#O��p�e��Pە�n�-xfϻ���fo{[y�/N� ��(p�����=����)(S���*+�l��vA���š�� �29�9���ꑂ�������%�n���#b�ґ$�{F.��>�`'��%��R*���ի�(���W&�͒T�Q.px��#����Xt�Y1�{i[Y�_�B|Z$�b�����!b�O�CJ�!��L��9s�FH@X��S�:�{�e�#]����_�Č��,�)��D�N���\�S�w��\eч��U/Ö�B��\�-��D��	��/��z�z�~xC�x�5�.�}���%��b�AL��x��W�*"�.���:�[�(I�����`m�^K��QC\,G�uH;�!q��c
���q�~����H]"�g��7�#�q�)�j,m�9D�#���=;�=��\�	�vT�D�*SС>^�߲t'�l�Մ��y�F�4K-_�����+������EK�JHy��#EUeR0v�q{�3�X�eM�Y- ��i���r�#�2K�&�r�4�T�;��Ou��-Tk�A�-0�)�+�l������Y	RY�Ɍ׃nf�Ulv���m�&g����<��ɲ� ��{Z�YTnS��4؊>� ь&2�DH�s�m��.�+kP9��3��c�LL˾��ϖ0�ݹ]g���9�G1�)Ekѣ�$V��=���!8�{ho��z_@m��tt��>u�h+Q�`�-|[Yy)y���>�;�(b-�dM~2�se��S��� ���}�D�u�O��ڻ�}"��,Wٱ�f|�