XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~��>í�R#6�H�ep�����WJ\j�Cm�������7>�PR'�֟��!����Ց���B%���D$�~�5����z��J��P��Bjd��+�P���9���5���}�����nn1���W񚧨nz�t�`}p�3��=�����Y����:����9M?��j��3�&c>9���*oC�ȱ���/���9�*Y�-R�г�f3��!E��[��W�|(����5�D��T����qv�R!Ԅ� NO���}0͇PhD�'�.}j���,�Z �b-~�'�Ԭ>(�2�^n���ZJķX�n�{!=��P�O��x�jT�Ϳ����
����(���3�^AN���MV�*�ӠqAs_��g|كs߂t�b�Ѥ�� N�j�����T§ESͩÉ���� ؉�ݫyz���^��B��d۝�q����A�%Ѷu�5�G`p|�8X����ы�ݙ�o�)��Jrg����c*UP���_�����	#�{-L���3��@2�[=��G��'1�_���E9u�w��EN�ƭ�$��IV��[��J�x����2����Ru&�CALs�8]Edn_������5��6� 2�fQ�?�<I�.5���n���ޑ�H���Z5�h8q�
p3�"6�� ��gX�#<� �v{j�
�o���B�U�J=�܍v��FX���xx��(n���Ru�S�y��r�[B]4I@aA=�
!�0��l�6����ԝ�]A������Q��]�1��cu��XlxVHYEB    7783     c00���h&�,��+*~��n�����$@����hV��B�|Ly&���8G�a1��q�S���ā�Ǎ�f�56B3��{I�+\21�V��$�Z9͈�����e��Md-�m0ɋh�=�n�u�n 8��r>R��G���G��ez��×�@SM���w���B��nV��vrfz��O.�A��M�Lb�+{��n����v͔�Wv��.*	|)�̝`��V�V�HcQo���M���⏊9����]M�y��G4��l1�M��	� O7[�@x�)�F� :o}sf[טa�1�^O�UG��x�^1R ���N�#ۗOn[�R�n�|�6�N���#a��1�#��4?�3��'m�������uG��f�����܊."��g�J�{�ԭ4~�	��+-�c/�{��ʦL�Ր�\���xJ��ʆ��`с��"J���X�_<N��-�P}�L,�6���ޙ�3�H���������߳2��0־�1�
��T���>96���i��O�$�;��W��(�g���-�AO8�u'��d����؃�I�a���`K�M��T�K�5��&�����/��C:��mr�}�7�����ڕn��,�^�_�9x�Ev�,@ڤ��I�=9FYj�	��2��m�3���eO:�� ^{�3l����'�������o�Ź��;>6���3���0̥�ݶό��um�|�Y�B��$;Hz�^(n�K��G��h�Bx#4k�]0JR��jL�ߎO��u�k�}[Gb:���փ�wH�(rW���|��
�IZ�)�$��)�䈨��̺�,�w(��$</���Uq��^�x�[�h��h��t�9=���H02���r	���Ց;��RS�1eIJb�$M$�֚r�l��õ�]2S)��-���N0����0�6KK H�Ų'j�I�2��E�=��r��.�3�릢���;�9Y8G>l�l$�����&��b��X��Ƚ���9P���q�x9L�P���[�+����^"��������9��Wn�Y����0*[ec 3_�^���w[�$�5+'��)�VȔ�*c��K��|��"os��P�i���:��U��C��r���٥H�jA���j^�xx��<���C��ĕv�"���a��=��ڒ�?�+�g`�MG$qD�e"�y="9Va����2Ϟ6]�?��	&!��U����0���d�s!?$ ��G����l�#�U|�j��)��K�Ы�r��O*��c9��Ji�	`O����Nd	����=T��$.��1�|���UCE)��� _?�R9�&,�h����Ξ����H��$q�!��`�,��DA�IcS����-�/(�{-F*����{� ���~ov:��Gw���.����|�����5���� 삄��8'O*������75ݵ:��XAd�'�[H6�[i>�Cz��9w��fX�����-RA�\~��[��g����`tz#����P�j�
j��������ҀBmY�~O�݃���U�?�ZsѬD񩦳��zCr��f';�N�=k�V�����w	��h�F��~���������^`t����K���8�uF ��'�%�:�3S�]Ke�ׂ��5}Km��GU�zF>�5�LȕtV�g�\R���+,�t�߾�(3������f��\�s�ϐ��zn�ð�]O�"6��d�5L�4��Փ��w��,mVD?>��և�_2�+�0%Z����ѿ؄D}�Ffj�a��6km-��������wY3GbI��ϑ���Z>�)e"*�������O�����j��7t�5Y��6*��rq%ٜT*�0�R��~�^E:%O�2X"���Љ��1�"��ɭ�J�D�o�	~
�[�m����h�7�*�J��~�?�9v���l��bO}D���"�ø¯���|S�W�3/�R0�k���E��,(+���6_�c�x��f��LV�1���W��%���FCð{:��d�,��E�y����ݼ=�7����y�:B{0�'tѳ GP:u���?:7��u7M�s�_��+�?�����J��g
�$�YB�T�亳x���U�٘ ���g&#���h ���� ���0�O�Ԭ:���x�Ah���0b��Zx�}����,��nNG�42�A����T�fr޼���'�-��8�|����/|��okB%t�7v+|���ùYԑX4� !5�RJ.�{L�3먍7=�k�O�?���F'$�,���gy0�?r;��%Iy�`�(N�ɕm9�����I���nW��a Z�;��X\����Z������G�Mo�_�'�_ն �=�����љ�=� q�Q����!M����u�d�^)���{2'�뢈���>��4��l**�^��Q��F'!�i�����+}W-1�L��&H�'���ڮ�i鰨��@�C�8c!��_NC(�[��a|�{nR���6���<,�1UŘ@�݃Hd�8�{�mYmZ��Z�$u�\���8�S6M_����{���H�~}h��-R�B��S$�h����9tҏ�v�����So+�
�ڻ@��{<Y�؛��m`��v=-��e�6���Z��x�j�@��\[�y�Ι��.�8֍���'���G�l< `XϚ#TU���]����fe��ӆ��fK��j<$,���F�T�	F���'`��џ�Uml������k�a߷*���u�i�R7b��'�7�Z�`�� �L��ڽ�Ԓm��܋���Z�	�̼�'M_���ࣂ�ĸ^,{k��.��N�@�&��ˏf���g�oY4����ٲmÚ�Q'P��-��a_�Rl���ʪB^o{���;J�o���6�I�}��������,��@^��8�:����䡒�<v��ۨn��5�no/��[�xD<\c%�8��#�h�v��O"�8&�����j[8�2���Z8�N���G��g�xBj<�	;�9Y�?[����$Fq�J�J�@����i�E����F�