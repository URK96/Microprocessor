XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%z�6��`+Hu�ݓu�'�<5�Ln]�j�P��T�_���ax���*<l/���`/��s�&�R� P��T ���z���G��M��B�*��IiI����%��73R��&@.t�~�$������%҉�3\��}6Q���bb��VGR��3��ď����ȉ�}��嚐��W. $�"�\��5+�7p����@fG�RV�H�IG)�4��ꚩ���!�D�>Fy���u�L�_%fc���O#������=�"� �
��KF'��ZF;==eM�'3������=��=�ʚ��>���ȏ����D?�ܘ�I� �Zt�eC`����2��B��sn&|Ϻ;i�Y0�!���PE�N�����sYC��W����9&�g��
_��r����N��K�H-��3��71�D���k�$��܍�@��t�ZG=.�!��0>�0���w����F�^5��M��Fή_���Q�YN=?����\qFy��p:��J��vZԭ�|���u�KQ�w/�����9y�*�d�Pu!�&����)g��/��,Z��?h�m�y���閈x؛�`�4�E�����	o���4�W61���|���f���f4��t��/��V��XM2��0"���_h2|8��|V쫝�K�ih9� �d����o�a��r01����
Z���	�|�[�1d����I�B�Bg�+�iX��������N�M�\T��#a�[��N��Q!!�>�v��&8�,'�c��ޣ?���W�%�?XlxVHYEB    4b0c     d60���E��*lS����z�Jp�K�)8(����b��V���ި�S��[Z��I��v!���:���#�O��s��kuB���r�3��P�i6W�P�%!7"���7���S4Nb�J
�~��s�f�!c�@{6$�� �i4���K�d�(��t�:���LR+��,n�K�n>3>��ɡ�H����E�-lPم&yN���eo�z��AԠ�g���s<��r�zI�u��&�>0�(<��vo���������R�5?n?��%�v���Y�������L�uן8��Bg��>aAA�w���%�b��D���(�����@�u>�׉�C�$�����rq��'�n��|O��=3J���.+ٮ1cC `�u*f�p�{��s�65FOֹ��.*����|���A0��QF�PB�C�{6()yZ{�3K�wT��`�n\��<��/_�;酃5�?�4�%�Y�,s�B��=UPiZ�C̒��b��?h���\Lu��j�2ZP{܈�&�1k�g|
 ���������^����哎��Y��a��=d�\R��`^�0������
[��\���SN󥚽�r��Mv�m>�i� lZ��W�h��	�3U������l�4v�#�i����>�r��ʠB��/�Qo/˖`���S#���.��gڝyV�e�4JAߪ�=��QIjx�0�Y!+���K�S<�������5B�(Y�= ������
$�g��<V�k����+c������ma�>| c(��sy�X��~VHC�o�el�i��@~��0�O?^�gn��m���`�����׳��3ܚ�����~����"���L��۟��"3A.���sNȘ{+U�x����������.���������	�n�`9F����ƶbh���'5�Dl����$_� +�{Z�B�O�:����#���D��Ca�����nȘ���,4,�=;��^;'�?_f�$%��1�e������W�g!D��=�.���(W<��j^�O��,X�̾�y:�����V�(��({o3QI����9�9*�P�8 �׼�y���9�Y���9���[V��}����6�M���DWqN`�+���|�A�̄{ˊ�{;�#��}�ǻ̛',p�o%���3���&Q��6*�n1
mJ���<�y8��e��Xg���!��/e����Ry~��i7=���*�}���hK�8n���#9�3�q�'�;���G�3Enwt���T0���J�=�����+UXk��&\�$�J� �����P��53/td�":R���q��CuJK
�}Y@���1�Jc��M�X����&�щ.��;�����y}�sk�k'���E���E���vًϨ��>@��ga�����:�7��	Ę�s��V3� HͶ�H0|[�mv4J2�xg�*�o;�s��<����VM�.^�?�Ua��w{NC�/j;aO�I��*��ʙ����i�fUx��U;"��f%��lE]`'�o3P�AV�U{�7��I��*��f=$"�x�H#5�WH`��5瓜�����e���Em�)���̨m`����6(�>.o�̫ۢ��|�u�l��)R�v�P�	�r#2H��h�Fh�q}�� �O��gAX��2
p&�JI`W����<��!>���Q��I���6O�H��j���k�,u�"�����H_��/�	�����[�Q=1� hG�jhRGe]�@�5� `��HC>7�^��z�|�T��Y?��g��?|�M2?��i�?�B)���2A���u���ӄ��k�`�����f�>k�{b�����8��
.�I�61�u��i��&�h3`���_j%�v	�ˠ�u/3P�p�Q׶�[���eb�5��:����4���=8n�8���H�;8����������,V<l�B��O��L	�Mj����n���(�挼��X��*�?c�6gc�~��_�H��5U
2>
��^KB��U{ `����+R��%�ù~^&�s/,��4��3Ki�ȴ�w��9�F����n�fĶ'���ND�^;�m�!��m��(�-vڣT�O�3�R%�3?�w[9�E"���R�p�kW�&em�=���#�,,T�?�a���>��!_�+�'�&%o���>ƠtW.�?x Ì�;C��r�w17�ح����BWwaS\� a;Y8��aV>~����))�~��lP����̱4)�0!T�;~]b|�<�o��W�83��nKQ�U��u���N�H����}|cp�s�9J\�2@Ю���]�����|Gӑ��^�A�̥�dZ��{�:<TP��%�l�=J��~U< �g����]̿f�|��#���DCj��GvXnޣ;q����0�%�L�5g#�ZôѺ�r�A�U�x�-4X_���%��/�	���T'2�0�WV2d�[�;hҹe4vM�C��k`(��I�����@� ()�`<7�Qڶ���n��WC�@��p�"x97-�Ry~���]�%���U�晻`ȵ;Қ=�?�E��li�!�N��g�����M8�J�(TQ��Z���5-�`T�x̡��i��!-��'�i�ɾ�m�b}e�0���F���%�>c�`�X�~z�,��F�vsjn�<vuX[>nQ5V���\4?�p���?��X����=N8v��|6E��*6q�S��d���泒�e�vC�I��!6OS+8����b��� X%� ��@8�6c( ���|S>�S����-�S��x���V
��ߖB��v��.�Eg��X���_y�9 l`��:c�B ��W�G�a�
^�r��b���������M_�<�>�7�,4���0 <��Y2�gk��L��X$G����D@X/��0�G�[��X�|}9T�^M�sF���J��vҾn��JMs��<�� �t�������EcU�(�V��f6ibJ���_�a[�u���5�-��3��Wc|\�$3���A���u�'Ac��ֱ5�e�����)N��QbY{�>]���*��͵[f/�7Qo�i�ZTc	I����-�x/4��	�Fp�����<��~����qN#��B)�I�9,����A�h"e��=B7a���R���ԙ�&O�����P'�y2JT���&�La�����:b{k�B����qQ�|�Z%V��Ȧ��:ױ�����Yn���<��by��:��p2%�{�Ϸ�� -�6�nS_�E����C��[�H�Z��a�# )x��sbz��iM*�2ϠY^J�	�_{nѕ�0J3�pQ�*� ��UZ�FS Pg�Xt���5���!�8����N&xI�$�F�kn��&�?�2=��:�U���tp�.u{t/b�H�E�����׳�Pԅ��5���3�����v(����-�