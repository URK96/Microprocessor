XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l�W��B�(J�ӵ�s��X3������!��e�7S�/ ]$���<�>��ʹ���̡	�
�8�Ie�p���s����Z���%EA�wK� �V��#}��vU���z��Dhߚ�����b��:F�2K�O�1@��{� ����@��4WQ���I��r�o�<N}|ܼ��kx���9WQ�Q˴O[��]��P���ˋ�
ƽY�%�8G�v��SQ3Oփd� S�^rƺ6$l�"
��#�J#�Jxz[���A6�?����ے5Ra~�i�\(�����Ƭw�|��ׂ��T�W�υ/��g�U���煱�u�-K>@g�$�K��P�L��
Sm�l�X��h��CEiQw�B�e�/E�[Zw�u�B�ġ;6(�^6�B�5||��S�Y��X�����]y
�4}��⡓D�9�a���)��"2M�=�雙��Dfb��4/]Zf�������:�x���]��y���5x�����s�ʉ�����j"P;/~t	lԞrPƄ�\�9s\��,�m�W�%�_���	�7Y�褈���mcs�����U�;e�^q��j3���̃QE8��J3�Y�}�������˙�%�����c:��v�u�yA������_0�Z�f��f7�;c��5д�#��Â����\�W��Y^�0�f}��A�&I�����&bUa�����<��eK�������tba�(��1!f���E��Cn���8 �����d΃�T��?�qXlxVHYEB    3248     930�x�%<�z��u�׻��F��C�LR��Usa2�$��n4<$c��t���|C��Wt\�w���ʹ��ZY��7b�Lʌ"PMy�G��b�*�k;Y�.= �A�E���3lo������ؤ�"��k�䥵t2��4[���u�ŎTT]poOL1�2��z�:U��]��T������s���s��#݆��B�gC�K�y�N���)��w�^�_��1F����ea?o�T����"�����.%�k�>o��c���hgh���Jn�r��Zv:�͖���>�������ƽҟ@��]�{����V�r�1Cl~��{$s�5�?n�h��"��+	"�!ށ����#��Q�=�hҴ_��?J]��0���I�fE���`�T9�`N��!MS�zh��ҳ��Q�{ U���.��Ć��!ٛ��w�ٺ)���iz�m*��c�6����^�Z�+#�񐣂tv�\�g����7����������{B�{�T�Q�1�'j�W#zA���X��}B�s��F����rq�Z���JX��ȡ��D&����o6���*���e�D����8o���	6�F������ecƣ���_�� KHD���h!*eS��Ћ��[e�q��T�'��F��q��������sɩ�7�qU��hN{`-�����O�
V
 ��1��������ߕq0�ǯb���&�uנ����y�"��а;�z���� }���C�[��@2��J�*�i��U����q҆L����ז!T�"#9��ݔ%O��a���V��c���XPw�y��C"Bc�F�2"5}� H�t�ps�-�	��e���*�����8~�2�7]���`;ަ$;ܠ�nⷷ}��b�p��(��ϖ��gqLY���0�U��#�������'\�+���I��#A����y���i^�X�����Q��Έ�6��)�FEӆ��ۋsu}>��'�Z�3X�+Q{X��\�6�����eȰD��D%Ԋ�6*�Y�d�
5IR�7	����k$�W}��l
w�_j/q[E�����d�1���̓^�q�-B#�dC�z���C�λވ$�1C���y.3��$��q�gl)Y�XP�
c5�s ��e�#��"cz[q��ь�R�M����۴ŧ��+0��R��~�@��q�;|9�'�Ӊ���H�NYq�$�U>�a�VL��}�
��ksr�d�����yZq����vnʇ4�_���d�s.KHԔ
y,kT�շ���Yنf��,?��tq��jj9���H��;w1À�՟3��<���z�'�D��=x��e;��k�����B�0J�Jv?Z6 ��,+��i�7�2������mn%��d,<x�/.-�S��-��#�b��(��V�V�s'h�@���=��`�-t�T�
�*�,ǟ�E4���v�����Yx��3ơ]M��K�(.��-��_���f7��#/��
+�k|RtSABD�)�,��n��5�\+�㵹--�7�әk4Y����"e��F�LG��`w�2 �� P�]����`:!@�}!C�k�ȹ����ca(�+I<��'T���d݇���H~�p5rʾc?��a�P&ٔR;��~o\�B;��-й�wE%�Ȱm/��,��e@���DMɀzPo�=tM�R��|���
�#A���C1`�����L��C������oD;�~'��O ��2�<Lx���E��-1�;�r�SV��r�byzQ)!��EW �����x&�u(fG��./蠻�B�|2�]z��:!��kJ�Aty�bY<<r���!DS9�B
'А�(K�Vei���������r��Cۿ���))	�!�j�w�^�r��~�����ZVX�6��ә�k����'RXyQ �@7����M����[UW��[0��=�ʴ�� n0a�n@:�B�Y�Gq�,��.����}��2� ����n�I��/�q������+��F�`�'*��gVs=.a}��V���ѳ3ӼMs���z���s�����Z�5{�d�l��#a��㱘���W��ڋk�x�em�Jn�|&a��g�7f����	H�ݐ��n�2w����0���Y,���(E�c�m�#�T��mD��z�"�o���U"�KS�@�ý%щ���6@��Eo��1��mZ��tP���La�Y�Ȩ~⁡�ܦ]���-ԃ_�*LN�{_�"�����&�(��ҙ@��I����S6k���u%��x�^I_���խ{��eRv�ƫb����	����%�����A���/��