XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C��!���WO?oK/�@�����շ���?��.�a�x�Gܛԝ�pUɜ�I�G	6��W�N�RM�S)�\^���S�H��|"sV����GZ�+�U4g����c�}�8��&p��	���E���@��j@���F�#���HI�N�	t�ψ�%#��ļVԏ�"B@���8j���B�����m�.+(LN�6�[ո�*����S��}նH�h�=�b��G:�{�5��_|��}hڈ���]�Ճ~C�BIдq8��>��_�>o`�N\�v�W��݈��UJ��M���X}}C;��zo�_Qabd�������C�@[�˜��w'���=����2����8IW��n�SU�Ѳ;�(�b �̜8���y�=��*��f�w<R�-ޓ�d�_>�E+����^B��������A�����0�͌
u�&��!Q�1�7��c�?J~�If�6�3�+@{�C���������3�-��h�A��� E�!���!���s���|wd���(s�k�g zX50]�@��<��9l����.u���� A��d+��͖�6d�x��/���V��H;D��&-G�%�]��T��y�������"�;��y�0ŋO��9���u��Ej=�࿔�E�9�=�0(ǟ�&=9��d�Ɯ3�̶��������c{�t"��aբM"b6���fA�;��}��GA2��}�N-_Ei� �qt�?rdK?�6M"PX�Ul��7PJV�ğ�GiXlxVHYEB    6d0a     be0����[�j���}���|��_l��Č�-�(�z!Ǽ@Ħ�E���,��З�D���<�!h�|gV�)��J+@��R��	�̠�J4ߤ*��IF7��ѝ�'��N`�����Z��Q{��c{'#X�+����Id�ƥ�+�>�Q� l�����2�\Jc�Oycz4*Lk�K6�<�mG�̓�G���vʳ���«N��D�O�G�b�d�e1��]a/f��M�&�(|:�Ǳ���Y8���wݥj;x0���W�P��~0�\fØNOݔ,�C$�c�`�""ɽ�ɘ��h�Ä�>O�mOӐ��r�d�o�^S��b���5��SD(��(`�q4[L��=:I�D�U����c�DZ;Q���;�E���C�������$�B�/�{v?���ca�T\J�c��rT� �sW(7nܼ�_�mW5�;���I{�������h�+r���"�%ŋIZ �S+�4T�x�����G^��d�YPJ�(�"ړ�1�iOIz,�����D�<
JʲϿJ-�7�
��{'8��C��r9mگ:�88�c����nz3��R���\���uP�}����Fd���Da;�ύ(����%����h�W���Ul�b�y���@dc�L��MWB��2�9��ٵB&I�}�1&���;�eT/W�������G��邧�S���`�����SՕ���Es6�.Ћ�=��׷O��DƟ�t����V��6?@AS:~Z쑊$��lg����f���T���PE@�VT�C��C�2Y뚱7Wt��;@�y��ǚ�<��}u�P�B$�o��|_P}�;��t���|�c-Ö��I���`��t箾L�Ƹ�.gUV�b 8R�bћ���;��K�]*�<��ˑ(��e,7K�9E��%.P��/ƥ���Z#9(�mn9vs �K;���b���#��؂0Z�Ԋ�j�ӳ��e�Һ&>��f:�D��<������ԇ��gїC'�?ML3(�w�����}���=��!�1]�a�U�WA>�����l��K��������`ޕ���q	�-�0�J!��(���G�¾.�)�Т �G:D�%`�h�C(��y�"5`>��n�� �%��? :���:�-��U;_��S� t�(����7$���R���W���;���D��q�C=�Bj����#M���Ld��O���`�|�&���$��Te輯?tEEfq�҃���-�#�\0Y5U���U ִ���B��b@���9��Bavm��c�FϪ���>��z]����a�&��;!����� $��'��z �y�/�����O�����W ���&_7�!st��}!�}�Ӓ-Z�V���ϼ � �V6<�-A�g]FH{FY��^�]����[r�ډ�[��aj�е����yl�
�y�k��gkڔ�W,�6c1�ht����=�Q��U8�Tw;a�v8\OҶ5s�Ԏ�av��e�<�W� ~4W��\�l��`�e�k�)Z�[���]}���C�	|X+< tkl�@�G���K�R�ȕ�зUG�`;P��)��~ �+�7�>h��I�za�h�%R�܆zb�.~�r\!�E��tZn�>�SW����P����\�b��Jm�U&A��F �j�&wYbaos�
�e�=fﰿ<&��Kc����\Ʉw�7�\�(��J�',���k�������V�1�����(}�R>d'��#�!���0�E���i�;Ōu�6�¤o�l�;W��PrG���M-xPՕm/��67�����*��8�ś����D��3Ʀan��u�1Ť�ˤ�sS+���Ik	"����d��.!C�8Q$�����^�7K��ݻ�>��7D�ta�5
2<rܹ&�HV�_�a/.��u�lG���'j2���"�3(Q��7���͐
I9Q�+�`�M��-� ��sn�!9�R��׉�aa�#�֗��?�V�f%�GEn>֝{ڿɯ+7���%nV��,͗��F�{��(¤udY�E�1��!�k=ʦZ�grl絔�� ��?8��VA_��{����H�^>����Seڸ�c��!�/K���!�:�O�Z�R=��E���{D��M�TO =m��M��d53G�1h��ˮ���h��L���S�.fMt.��?R�XIIB2_��� v�zF�~��q�����^��Q�NC���ĩ���@�vx�����`G�A>����ӍҪ���ZcG$��ǯL����%�( BW:����&d�ӊ�p�-����e&õw_�;��\��)Mv�������cb��D���FmI�}����������+�|��v�2��"����iA!p�L2��Y��v�}��	���ʈ���k��e��̄|h��z��%eO~=���ܓ�W�3(?���h��jYi*Y�)�P�?�?�_�l��$����~f<�=+(�oH�א��I�m��b6��i}hT�7�d#+O������itu�ѮP�y?s=h~�mw;He�ro'��R�K| v��j펋W���ۘE8�^�omL�YB����ى)�X@��� ����ݛ�,^��3R)%��6�(�s�*�k,.M�ba�N7�ٜoE˖M�b�����lY��F�{�VG�H��[?�^�xlo�1������%�W�^��$��B1ģ�>��f�C����y��5�J�H_��?�x���ĥF�`��Q+K�e���g�3��:�w��~��TO0���eNe	����Cr��(@R�̃P^B�Q�뿈���QPJ@Sg�8�\l@-É8����f��UNh������5���������|s-��� ��L9�&P�g��ߦUȆ���E���_,�o��|�[�+�K#^\��"��)�t)ņX;��#�`6��^8��Q~��� t̴��R9��S.} !i�sl��k��