XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G5v1!]�O����yw._=�z�6]�,��K����d�$פ�Y*%����6��	�'kdCǷQ�˖xB���2��8��&�I����(eR�G6UB�}o�"��:��wF � b+�g:p�o��F�(�������ܕA� ��S��/��f��Z6��������1Pa�eh�*�L�7��MMr��,+Ś_��0���'�f^��t`fh���Zʷ��0:�Z_z�غ Ъ���!�ش�����m^lR��1ˠ<4���6r!��\X�ᝮ��;u��y/��ϔ����2I�-�������@Zޭ�/Kx3\|��dϟ0���-�ܘlLT�r�.���g��@R�q�̈���H ����	�� �L�S7\���5%f�w��J�p�sK?����_��.�cq��2G���9H���\��@�N��Gci!�lov��b.z�.�������#3bl�PÐ���H����d�����@g}��������_��_��l�߻>z�O#�!�3���'h���v�j���~o�.bD{���s�0l���O����O�&��Ɯ�s�YFN��ɡLRm���SI9�&���� ��X���N��%�Ok̒p`L�{�cfv��Ϫ�|����گ���Y�u5esHjֿf��n1�����#�l�=&����!�8ۇ%�Q� �W:~�ˋu��hT2�mN��_�9�.tM{T
����3iz'�(�05{�>�r�J�,��{�@f�x/aXlxVHYEB    165c     400�eO��:���F�Ykk(V ߶�����l�ɛRl{@�$�c�]c0�Y�q>}�C��xd��)N��;�3s`�����z,W*b�w0�[רtY�W ����_�2�ժ8�-}P$�ޑ��l�`9
WHw;YdWw=h��d��'e�	��e��T��4�ںթM~?s�8�/�n��,�"NIV��1��`Xd��C`j*�Y�/�P����Z3����O��ߙ�A�&��������cҷ�VLݦvs�Xx)��\��x���n�5#3Ui�X��'��i7�)͸�Q�}H�V8Q� �W�"�T8���2v1�����+xUo!p���E��(ۖU���Y�	<���J���&��]|��&{���3���C���Eq�+� <yF8*<���Z�?t��ߠ$y��3�����S��4�)��v��F���}�9��^��5�w ,�[�-l��i�6V?K]� ��J�ȣ�7�Ў�7Q;��03Y{��A�b�Ln0*Fe�a��W3V�}��&@A��R�ޡ�'k�����N��>�*?Y���&��5����b>�B<�@&A#}t_R`J�DnS�I��E�f[�E��sb�F�,I��u�4���ī't�f�m�Lo�~�,�D�ؕ�(Uen#4��Mz&�������"YK���ʝiO������6DL	;Ax ]e��iU͡�cB4f��Y.k�Hh�[2)qH�XW���G��+.W�� ��C���~���.��E?��bW���([y�Pz��^I-U�˯<PD�>�a����+X��~bQ��P�'��31�
�>�^�@~��^g�G�?7s�R~�̵ܼ�'(�E>Ja9���QyN��%�襛���F�tgՏO�c�?p�&�D�z�AaP�&��PU��N�a�H4��K���-ڲ.�	���50֑8z��Ө���ѿ�Qb;݇Z��k��v[uI�w�f1�4[~�������j��T���|���o�D�)R�uF�{�^��y(��e!�)���