XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���\=� �,'��_F@tq��O�ێɁ�S��U ��.qZ3��M�V�b-�5�tn�$���=�����aS�d�8\�F�S^]��"�%����>QZꖡBK��6|G7	j-b�1�s��1S���ǐ��6�9����b��{���w����� �:U]P�%F>�#-���I�,j1,���E��ȿ�O�n�-� 9Y&鏃s��z�(U���6��3L�]�X#M���w��^!u�o>ٹ<���L�U ]֕����0���n1�-*�q����>Lfg��`��C@Q��IX�z΅���b�n��;�"߰� �MG��A6+ʀ�#R��n���#�6b��b����)d��(�+��PX�Q�P�cs�~}��V�i���Xy�6��3�o�ȕ\|rٔ[.��I�y�/�c�����>�f���jC��M�ジpR��9γ���/dIeYN,��m��F�6��Z
��(T�|X^D�
�o�JpG	ZQ3�Ȍ���@W-]�>�<)ے�ywTQ�s�l�����y�չժ<�`Ռ���6�>����(e�@��Q?��3��͋9Y$�53XD�P�{���=�ַ���SIaC�?�����ԮoZFG�����@!�����!M{�u_�|"��-1�$��;9�4;��nz�����:|qn�p�6�"�9S�����I�I�>���!�?��>���C��KP=q�-sJi��	GG�C��_6�,Y�:�kш�H�+�[�muXlxVHYEB    216e     8e0R�I�,ӫv#�>8�%.M�A��f��K�S���V�ӕ���SɟP�R�U!�o�F����r�|R��ާHCC��#qk=�[G��g�h�#�i�'�W���SG�O$W@�%��ċ56i;�4�7Jh)g�1���x����(���?P;A��N��y�Z��ə����*��N`���b�ҖH3�Y��[~���)顳��" �hbS�t�6��K��W[/Ӯ��]LK1�2���cxB�@��X���g�b-�m3~}�?�����B�1�H	J��U�f�N;���x��~�n 9&�4j���]���"aMXd^�����2#Y��H�#��6&�j�e�ݴv�=���P29��x�[Im+Ԟ�>�U�2)%`�=rkG��m�����T�X�my8��C/QC �Z�er3��̥���1��s�����t�_���Fg�zB�&z�(�_br�ez�-�Aq3������U60�qs�j�f��c�E�bh ��?�S�ԑL�g�է����ͼ+� Mi���"G���2��ttV�v[�	U��023��;�����{a��!�p.������ǘUc���!6ȏA�ߵ-%.Q�����k_A^���7����ڀX%*`�JI��>G0�Uq:<�+)O!k��h����ae��D�!�pDf{⾴G#� �J���X��;���.��F����u�r�UsC���!�s���_q�g�j�9Tp��w��o_h�f(kpQP��}��q��Dp0.M�h?�s&r��..1TA�x��)����Ȟ#���rl�9�|ȹ��
��z�C���i��eG��,*Z��Z�]��PP�H��x.�:�a-�\���V�A�|4ڢ� fb��������z�H�x�]��A�Y�ƙ`��$-»���8�4���"����;�:U.bd��l�h�=|�5��ǧ�G�:�PX"B0_�^%.Q�*̾�����S�"�� ����@>[�f۬�1� (���J��	��dO�
+KYQT�J���T�,��aGM�zl���oo��ˏ=%WS�׭{#�!�['��\��M�@C��f�9�XrO59B
���^əG�mɇx������e�\��s��sA��uʩ�ڑ�唌����Ò4u�WP>�y@������L �b���<	��>
!*Yi-���âG�����d�!����q���y�����>d�-(}�%I 58����]�p�%7�aܛ��Fh�+E�U>.���2c�c+��K����JCI�����2:̱1QfU�߈b�����x�����'�������-9�|����{L�99����2��S����$��d���*�Ā1:��a���}��(��� 4 �	����O�Ÿ�\7P��E�MhJ���5e������fm4r��J��/�w���K���_2�q$[�h@o)A�����"��M��g��Zt���y�1!���g�ͣUZ����G��������Z�@�����QT%�@_?����=J+�I��@�M�O$�7y�q�E�^� ��Դ�W��r�qt"�&D�s�/w�'�g�?3��$�.��p�#�u�F˰�)j,�������c(�~y �$gkȸy� E��.`�M�dҮ֌[3'(5�|e��U�g���.^�?z?"���1�g��kk@���S]�N-������ۂZ+�D�r�5����9M*],��o�*��+~l{�ǖ���s. ��|�%�L82�f��2�1���91B���up��0��
hW�t��T��Q �pB|���',��~�����vV�������(U�V5�^$V����^h��+�+J���G�Z
 ��K1w��k�b��z���26��9�3(P��wS$��#��O5�y�$����c��E�!���^��%�]�>��[����q�T,�;��׆;6��iw�vG8�c�!!p�,�V*��INn�z��k#��ݸ0B�;G�+�&>�D6�� Ч���谱rWi�1�Ao�1���`�Y���n�yro_
��E�t�����6_ҕ�>{>�lȘ�gE��$N�OfW�,b��ֶ��Y��V�����E4<���wB��-����L�9C������^�~��Љ{r��:�^��ۤVwEAA������6���~��NJ���Y�V�u�͒�$��hy6!�
��p�8����nv�y�>�A�+N�x5�x&��6�+��(��M��d�7%"� �#