XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��gn���>���agt�Z�\��C��GtS�� 6`�Iuo��OU��j>�9�X�jQl�~p�ʡ��Gi�O��H�#�Ɉ�B�����A_/y�m�<6�BT�����Ϩ�<�*P.�p;�[�޺l�[xF@�~$�[�_8�,-��������n�P7��ܲ�EK5�RE���������N��뢝����d��I�?�����j���&��q4ˎ�d����"-5�ǱU�J��'87�gg�9@��&��	�e�A� q\m��j��#�k�Z�*�a�d@�xӄJ���M(�U���5��K5Z�߱MͰ�hѼ�>�<֧�s?r�%I9�~t�z5<UXW�	ǩ��r��m��F��I���f�/�.c���tn{5�5���2x�F6/^_8������N�ƒ`�"�ڌ���B��G��%�{���مpPcV�]S�.�7�,���0�7J.jH1�A3�jnW��W6�!�T) ^�3"�>���n��ӹA���+c���m��	�wgs�_z� ��R2wc���OL�:r��s��1�&��u��
9i�\� �C��B�gpiUb���	�TB	x�&Q�+�ɷ�i~d,Udsw}��z�H��ͩ����qB�
Ezi�}�*�̣n�Y��P_�@�Ҵ�Ӵ��SE��k:�9;H=73tA�ᄨJQ�=ˣK����[����N1�G��~�|���V�66t\�f�5��A=�2IX��X��)��g�ׅ��1XlxVHYEB    1d4f     7b02�=�H�B� @2�����Q����իV�3 9Oa�?��Ú:�.�^-�����'�L��,܌�_lZ�q�r�}KŞ�R�c������CٽrsB���?L�N����(�eQ�⿠�UY,�K0`�jx�RD�gQ��x�	QR~'q����c%{���V�Y���j����R@���eZ��Fp���-��XF"��c3b���. �"6i�j�ҏ��j�AO�R�^e�F���a�/��,p�Jc��͛Eg�����l��-2[zA�� �%.2��.Qӝ�ƍ���c��5;��O��Y[�uה�D��L�Tp�Od��h�P�VQ�<׋D�*N9���QG�Z��(��J?���}{�N�A�<1?�~���_H�����!�!��b0gֳ 䉙j��?sٮHP\�v�Z� �#d/�<��3r恀�ke4�-_f�>�"0�\0}̺r6|c(c@��Y��*U�G8�^}����Q�-�q'o����ypv77�*!^�W�~���&��� lnQi���e�����!ٌ�R��⼲�h�z0������hO�L7pG���EB�a��;#׼�R6Un7�6�P>��'���=���' ���X��Q�|�
�����'U�&~��1�3�0s*�R�p���ݩr�{��:5��>G����T�]�K(+�-�7��3\��W�<Ɋqv8���os�V��G���b$�O��R���v8{u�Yn�Y��bH�B%]�X��2s;?ia�B�A�.j%�h>�fBʶކ�k`��q� 8�[�v��KRs��8�/��nYuT�e�)�u�֔ޢ��,�\��2 6ȍ�p2�3G�������PA�ǕTfG
,�\I��FS�V,��OD�[>����q�U�8G�∬�N8���8���j=�W����̞]~�3����/IT�4����s��'�L)8��s>�����x^���kG��oT"Z�+;0���{1�9���<?I�!�-:�}�X}�	ׇm�.D���-�8'VȄ���D�YH�h�!�E̇��Ŕ��}9D�uV�L<��Z�[�̱�����T��3�F���xGHD5�e��X��+M����"��.̤����R��[=��Z����:HkA.��Ysf���}8<�W�&�7�~�*�aMJx}&�]!����U񂲅Xk�_nI�ܯ~Ⱦ��l[Nee+�z���dm��
��F����#Q�y���5�\��u�,�L��uԶ������1gu������H�S�:<��b%�&�vQf~�ȣwe���X�T�1O��㌚����V��J@X#��e�5�=ͻ9�ZK9��F��eKͱ��')�K���#Q�R�<Gn�B����=���J��/1�f؀���Y��C�xxY�a�,߸���,"N��������N'N��YViS�� �#��v*�RRd��Р=�Y��Y�ȡ�i���~�tַ���{(�C�T��3F:��kt5���,%}o8��r����Q�.XZ� ԟ���{;G�j�[��"U�ܚ�դf)1��f�Ѭ턷��m4�[B_�������/W� m5���	�1��F�b��Es���l.�>�;_/�O�+��J�S�o��	a�����*��"4��Zj+�#e�R���j�J<oO'�*P��Y��\� P�s��M,��V���ZӣE���'9���t5W���
�W�MY">��9�M�@iC(O6�.��a����,��hS�X6�M���<b����X4v<cs�@� E�C_�
�#� �'��e,�n�$�u:U�;'I��n�m	n��+2�y�QN���O�>��|���>ɣr�ϒ��n�]A��Z���#� ������-=�NS~�}��u;���S_��C�o��(YU=F�8E� ���)�I|