XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3e�$�����܋�i��!HcN]��� f�O.�;ZxB��q��Ґ�������<��؊�y�-s��Y{>��'JtX����;��QyL�cU����[�G�@�u?����������?wb����T��~l�層AW�v#2��_5#'���ݗE�ll�2�cM�Ν޼)Q�VQj�>Sʞ��Q�I��u �������r%Ƙ�<��k�_�o�h�����᮫)� KQy�N�mP���m��TT߄~jhҭ�#�m��a��A0wt5.;Gw�����Ng�-_�/�~�:.�rL$�t�
���ҬjLÈvޙ��nψ,%He�v䄋"��xj�aξ���{T��c��#�ū�/2�����Pg�.f֒�Z3�^�)�o���lq$n��l>|
5��Q
��4	 �Z|����$OԵH�$�:I�U�[3U���d=�ݿ.�~��"_����ᖒH8q�OQ'xuY2�d�B�qME�ze��!H�1M�'�h	��a}Fe51������>���E"��	Ȫ�F�(ڱ�M�^�v��߉H������&6O1NRpw�]4�,*#��P5ُ�i���!ي�����	5�q���0��z�
�(���Hy�����
����H�Yb���b�)eN�)�{J�Q{�Z��Z:���"�l�Tx��܈%~hu��4|Y8�a�oͥ�^����@��jz�n���!�M��l7lG�t�L��C�uf
* 4f������ڇ�?��@��?�����UXlxVHYEB    3c8e     900�R�WL��UT	e|v�rH ���ix�{�3�0a�Ӫ���;��k�4��νK�� ��4�l�������J�#S��?9(����v =�S�<�h*�Sr�h=�N��>H��J�����ė��eVy��>\/GZ��g�;ze�2:�GB��,�"&��}�2~E�s�z[��?"�_L��A�F�́�'&�b�����g�-� �.�̷&9y��Ѻ�����(aѱ� ܭDJZv�3B{�?0�a�0#������z����U�_�ϴ�OG��U��P��1g�e�݊��HQ�=�4�����"�Z�b�O�$�Px���wX�1ц\m�a �V�����ȹ��{�5I�_��B� f�e]��S��#�����
]W�}薲��x���T/��Ӕ��ыJ=!e������T��$�ϫܻ_��|���9���F]��#`���i�����C��
�:��x�[ec��ק�˚�V�-M��¦�3�����y43��/�g:!���� v-�6?(������
gIXz���J9Y �ط��yYR:B�Qu��T��'9G��
c&*�a��[-�m��ɜhXwa#/x�\h��X���B!��:T|������3~,(��q*��Kݡ_߳��9�ۖr�h�;y�F�4�wH����g���[M��v��'��%���w���Ƞj��3��T	Re(��� ��n��gA^�<�*���,�nl�$M��P�,w�p-��(&:�%G���L��.�������H|���'��M�)k)u�L�dn��B�����-�D�n���$�"�����S����]�t�z����#[��̪���3	(�����"3�{����gH��U�0�6���[>� 6����"�U|ʨ�:�eC�J)q"����O�+�}��
F��g����E����$�S�����Gv�����p}Z#�j\��o+�;�'��v;�TƍP�=�m�
n��}�����%5F�݇]

�G:�m���J�����̶\��$���-g�Q���VO�6@��I.���6�a��n� ����dM�_�^4��r�s��]2��y�ZUE	��$r8�;��π���kU.ݢ�}l��nx!��I=�x$x��C������V��C��I�XPu�J�yT��q�G���r����Ҍ�j?�@����5���M�aq$�褶�@(��L��9_��TJ 6�v8\�~`M�[�Y�+xШ���hG�=�������	��=�z�����T���͸i����P���l����	�4ul�/�VO�鐰�N��F�m����Cʞܖ���7G��C`���Y�D��;�:��G���	��~����[�	��}�*x�*2I�`�uO�ڋ}/�s�(G�O�[�0<�0�K�^7�8�0���K���#�-y�N���1kF*/D��Qs�� ��A�v�cIm�ROK�--�V���׆�ѷ�a�ܡ��@mL<����,���R�����BaLT�N>$&�r���^ZP����I�11.IYι%�:�A���O�����~Tg�!�hS�(/�v���Njqeo{�CBW��e%f/�[�����`��͝����v^��b����]�V)��jK���o�d������W�8�v�K�lE���7�I`KhpƔOn6���)xՎ�'|����9Y|A?5&?���"�ʆb�������xm1>���Tm�
�L�d�<��EO��{LD��sN����Zb
c��<]k�LZe��S�8�,�m::ᢣ�XUۃ����q�z���3�
q��́fUye�2\��F��'*�?!&0R�ݰre����xܵ����~R��J7��گBlP{n|_Y�Q�U�@\L�W�e�B�#0a%b�7����נ}|�0J�	��͠%�C?��U���s���3��k�k�T�I�h�&�6g�'^�ʠ�a��c�X�߳�ٵv�/-��.#�m�!V��C��?9\pcX�?y�)>�s]w�R.�8�ĺ�b[�V#`F��V�U���`^���tR�hc��լ�qJ�������4�^u�p�9W�"�A��A��p>��<vc|�P��"��������<E-*o�s�������%��IZ�25O����r��(��u";.꺗iԏ��Q�%���ι뤏,��VI)��&~�x��s���8Ѭ��T�[��{��>UL*�tj�Q��kzP�Qp���y}b���,�an�1�������