XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��N��z5��.%�U��1��Q�!����t3�q@��Y�DP�3���؂�)�{�&c]d�\���ᔤ�y�<���55G�/9{�ҋ��K;��wBK���~�e��굀���<����	�LlR��8OyBH�ޟ���=�OX�Vb�>f����ȣJ���j7�v�4�e��kH�#)�[�C������-�x�Zp�H��,4���������5P�\�@�u�**[��嚰��y�JI(e/��_ۙMx�����g%��.;����xC���.4�)x�2��T��E�ڮ�;����Z�̈́�^�+W�;�e�l}\��uټ�_�$}�>t�G������K��SO�+�������tD$�7�م�GZ��SVޔ'4y���\{���.{DiM�!��i�U���,p��T�aO�;f�q�<b��>��jڤnf^���_�uQ����&`B�l|M@�{�a�VM�H�.�V��<�K�u>�-_PD���
>p+���Ff�t@��kL������\���O�<��Û��}����P"e�BQ|��(�T��ǿ&��`�wҧ����/1?M���.����� �@ב��7�2�}��ܱ
��A�����UeB;wv�'B6�}�xX����W��#i.$7f�j(T!R��d�C���V��Czǉej����t��ֲ���@��Op��\V��:�oi d�&G�t�՟����o�p�����7�C�ѷ4LѰ�B��ay(|;XlxVHYEB    1620     6e0:������
y��r���@a�d -zMO/���9���o���^�K�[3ԔA��,��K�?�����������乭4ZH����$>������n'r�&��X>+M8���)�b	�X��K}�'gV���o��"t��o �������HNv/v:�N�W'�M���}Ny��l �o |��s��C�w�Nk��a�P�jN�ih<Z�>��Rw��eŊ��u�j�^�j�5��XL�H�S���'{�8XK����C�q]ˤ��lA�zD��t;�^µ��a����>$�L��o�?!39d!��<r>�	-��k�{�|m�H oF�FW N��YCd!񂜇����P(�Kb�	UXd��]V�$�e�����G}:A[�&�:x���9V��j<�8
[��^�@������ɐ8`��I��`:�����jjl��P�.f?"zv7��8�ѰԾ�ȶ�/���<\.H/������.�q ���!vxt�u.�f?�&9��dD�'S�sO�,ȕ�/q��>:/�t���OEb����ĶFv�6����_4�D�����-m��m��I�'�$�����*�������\���h������SF����^
jH��C�ZP���2"N�M���ɢ���+���0{*�0�a��l.#���x��I����$r�!���-����d/�A��Z�%F���a��Ѽ-KA;6��U����ZqO펒_�~��$1G�����q
�d���Z
%��������+'>K�B����p�R�)��­�N)����-�̪��X2^2��gL��{N�i4�E����O��l�]�TH��������Q��c�uߓ�����Uh��Q��!߯���l��
	�I �K����i�^�q{�O�/hP��$ ���j�Jv��w��:�[��fK>c���jK�4#-���9��#
*���;d �q_��2מ���V '���$��C�7mr�����6�ݤ�J�W��.��"�ccԵ�z.��K�H}W�9�U�M �o�|F��k�#�W�w�m�*��D��@�6B�t�V\MV3Sz/����^yw�
n0�Y=�QG.�0�E�f(��Z_��y�w�8�4[��$DV�G(�j@s��6�0�A��ϝ�t�x#\Z�&�0��fy"�5��$N�h�y׬�	wI| 	��yr���l�zl�\:�h�����>�q\���`�&MNC�G9�	������Oq��hڱ�9��h9)t"�� +�@����7�tӠ�/�� -gM	Hê	�K�:~;P�F�?&R&���m&�C��\{�Z�%��K?�v�Q��-�"ꃾx�G�9�:nx6����NLZ��4�Ub.NR7$8"�2�+�4��F9J�1H����e)��E�/�2G�!�(��.�vS�7���W�����̺�Y_��7��^�{щW,��ܡ���˪��C-T���sT7@-'t��y�����?^�~8�8�>+��t}��ůw�����^�	n� �1�BQ�.N�Ĺdh�T}��m��T��D���ÛB�I��K�^֌oy�U����aG�X�&�3Yb�3�(>��5��J%]��O��z�:`�]Ih$�f�	��}��sɚ��fMv�ǝ1|2�����@��(ű�):��c�L굔���M[��M��D��I��V�A���� �� %K^�׬$�1���AN��~f-�p�}��¬��40tA�nJ���4