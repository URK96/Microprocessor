XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���� Q��nb	�Ϝ6�*1�w�cO�y%��Jq��'i�}�o���a�����i_��kڜ�f��(%0l��]�ީ:kL�Y�����T��s]n��Pۨ�_ub�o�U \������Vё����AENNNJݱ����:���a�9�=z!��K�mtU����sJ��Nv����s����>T�%w��1V�u��<b��Iz禬�h�9q>��}Gz}24nN�ޥ@u����#��z6h�R�������{ ��8&'�'4��ogs(jL����n2�rъ��'�����1�4Bt��],�_���;,���H�J(`*�;+*���&����t�x�9*X������||�v�fZ�;�����+3�L1���!�|A�@A�;ρ0��[�OS���A�%�������ȥ�����Ht��N��eX�����\�38����K`�b�*�3,;�����B��`�%�&�)��ѩ�t��-G�&(_CX`�cK1G.���U��	�yo�Y�*�e&�����,�����N�1JQ�+cYԶ��L0����J��?�3�����3�cڋ	�1
pY}��ĚE��Yjߩ�#t�q�:��'{FK(3�L��,_k�����t��]ѝx��;��
cB��R!�K��Yܶq�'-��(�"Y2ռ��E�sQL]����p2Y�A�H'�Ws��M�aV����+w���i��2� P��)�0w��3�{.eϲ�a������8.XlxVHYEB    1c48     560x^*��;U���t���X+Y]	wsL3����	�2���m:�F����Lk�����{#���f�Dl3'_�w���k����m���a����;Z���Ǝ��9�����[�ݽEZg<Q��*\��V��1f�r��݉�X���ꨕs�s�挾�( f�b��4'������\gq���ֺ/�/MKO�nQ���^���p}QyȮ����`=h�YJ���[?�sm+�����/�_o�)��4�=�PNݑ�#�C�Ϲ'�.�jXI�B]���j�}��lӖ��_�G�m��̀�ž[�q����r-��
�Ơ1�4�W)XT��L�+�r*�W��K�r5TA���}�F#1�B�s)B`�Zq����*��٭H$T�:��.+�����k�a�3������k��$hj��C��=dؓ! �G)�mRa�5G0�E��k(�J'��v��t�)����K'��x�UMX���>fe��e~����e�L��s���AC����l�,����~��ȼ����9R���aKc��������rG��δ���P��/��16����G�,DJ�ߦ9���B�wLg`�%fz�#��Ƭn�{���Q��7IY z��F�o��^2�hhf�UQ蘥�W)�_�&z� ���p���~��s�M��i�dw����*x�
**�:f���fJ���]����̌&�G�sȩg3t���ST����2���2Ĩh�w�mn���WA٤� �^�����Ye���o}X�)_�F�cg�ۀt���P����Ѱ�#Ŝ�l��� �Ӱ#���q�L�p���U��#ƫ���Kuk�8f�e��Ҡ�� �� a���W�*�G�/k,�bZ!����[W��^N���ƃT���G�� �+�HT�O��5�6�W�/�����ն,���ac���;��ģ��,����o��>�f�1 K�(��~��6���P��;-)ʵfo���Ǯ/�C��>�2ǥ`�� ®�A��nsv��GK���-~�ՅG$Ӓ�4'-=Se�I��Щ��=�o��u�������d��d/~��vRo���N�P6�����Cl��Z�	ZC2U/,
�ʪj�����":�˚1eZ.QJpZ܈����.�0���kv�Z����:������p����}�۹��9x��d)���4XJtz_�8�~s�%�M�Y�n"q^��3]ä�����X���C�=g��t����NvG�[}����%�zdZɏ�qK�J��N�7Tb�H`�nU,����	w�{8g�.��O~ʆF���CJ�Kd�p(��w�QqM��Il�\��PEC����L��|8:^US]i