XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z�
���9C/_���Q*@y9F��2���ol�{zF�F @,/�Vp���T�3:��(�gL���m)f�nU�z:	�8�7;�C��=����(0��L���M�q�4«$M��+y�F_����].�q%�΄@���B?��t�vZ�i��S~/~��G(�pk�֣�������x�:s��ć�V�����+<����2�}��{DBH�}���b+�aH�B�l������+u')G
m�*?<�_�.��S)�]��-��m��o.�+�t�HS^Nj^�$��7^���JZ���0�
�M^_)2�Jx��`���uq�ރ�DW��2B�he�)Q�_�0�J�e}��%�ɞ��@��S�q��2@^�Ga5D��ʃ�~6|�!W���M\�6���׉��[��ev_��b�?Ѳ���m`���HAgjR���RB@y#��+�ר|X�)P,��x�|�+����"��=��-�W��Ĩ@�Lj/T�z̋����{C]�;W6H���K"*rL�g���	 ��U0���4�b�+�hP���"9�wOm�!��ɍ�sl������o�*ĺ��w����֟>�`@��¢0��Utͤ]뮵�х�
�&Vh�}�˱f-8���H�U؛��<t���H��8��}7Mmy��rCr�.�m*�L �gW����B�w-:P9�(y!�Z�Ax/�%m���
�/b��f��E�(��+���;��/vJ��&�b��4�GR�{=Aӊ�$�R�dXlxVHYEB     a4b     3706F����S˓1Ov�� �2��$�N��A���V\�Q<|���]�+�ϵ���5�0+�#&�!�'*�!
��������""V��� }+_�}�5}1=ԍ�d��4�6I�Q/ݍ �3���?tp�Z_\5��կ�q�cK��F&��B��J��=OoS����	È��ű�އ�S��8�K�_���K1fc�u�\�OnI�a���GT��}
}f�����ۉ��9������v�>��L��B��	_f�f��z�c���3 ?f���E�a^�
�<�HY���ԣU�!pH��9-6��D�n$C��5��G`^#����p�SrtV0�b�һYc�'Q���|ڽ��Ӧ�FM�U�s��,�c��!P!4@��W����9�V~RQ����^pk`�f�Q��Q U��Q�����r���=7�w��	L7[��nP�Y�I�{�*P�HЈ�\X.<yk$�7ٹ� M�!0�kB⾶kVg3-B(�o��`������	�Le��Sf�b�Z�x��W�^�E�Am}Fh�S�ܵ�����k�����\a�h1;�|��W	f֮bb?w���E�d���DU&Ǡ�&����A��8�ݨ��5=$�dH $#h����f���"��R(Cl\�}�U���:�'�fhxQCS	�����\���bq�����M���*E_���$��CK��.�ҚDn-Rr"�I�Ԙ�j3�|�f�~r��(� :y�L��Zdv�9�`T3CGW�B:~��=<3��U$�#*������$zݑ���/O7yA_/)o!�9#�a$��N5�#�*4.���z��z��ජ��
+όL�	����]��}�\:/*ؐ��E��Z�(ߟe1��<
����P������K�8