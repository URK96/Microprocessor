XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���D	u�AZ�$���L8U�]zѣ�@�5,vjR�����VhZ,,�k��h�ݡ��dX�pc�}�
�4������f;����P�AJ�qL9E��`�&N��s�1�� �~ �jC���j��X�F;��|L{�6Q�$�\���Lg43"=�-��C0=x[r��g�T��z����$�1��t�ri���*�f����2�f�
G�V��wGv>�*�sH�2�~�CJ8�z�u\���L_Wt^�v,��l��Z��T��C�c�l����k��%��K�u��� ���*���mo^P�+$Sq٠���F��c"������T����4��F�O�i�AB���h_{/�<�!�*��m�>��,	\v�;�1v����f�������� ��_��=�K�����<&�+�������������h^�~�C~Y�q�'(�:ʨ��dQ��~�Ww���`�o,���P�Y�GQ����
f��yb�+�O0N�2�U��i4��vr��������&����������q�QBw���<ؒ�#�2�"���d�8�~��X�+U�+��D��8ܷnN�4�49Gi�����5�kҬ���g�6�D!����k��(3~q~�i��x�p�=�;�1����ц� e�/e���NB_��w��#�)�tc*��<�X��]���u��+�歎���f��=�ܼY���+�~i,�c<b�c6���J��ut5ӯ�J13|
XlxVHYEB    1491     490��d}�,x� .,���{��4M����[8��w�$,�2��xҚ�Bm��.�����_�{�k���c[���'Vuz"7��x4�?/���<�-��z9�5�����CܚM%]��z�Ul�1�����lvA��w��kR�A��o�V���i-~�$��jl��|
㵻�VX\����4F�s%Iz�8O_�O{�� ��Q
�/������є����S�v �V1�&�G�y?�:ygu��(�F����O]MX��0�F���q�F�E�[��Y����j��.�����uBD���擽�r�Y�;�ry���)֮1�?��AC:Ǖ���b� ��\�ܕ��m��7��I�ݝ�["8B@��̚S'�1X���N(��D�dK��1���I��R]�nXZ�ňVZ�>�2̍���Z
��_��w��]��7lٔA놦��)��R4֭�| =>#���a-x����(�4���kO�"����$��s�Os{/���%ɿ�2]�7宠J�U�燾�W\ZF<���BV�l�?�h���t���9�k�l���I|ۥ+��GOљ����_:J ���Ja�#k�r�o�]6x�zf���X�?S?�(�E���&s7bzF�h��;�e�쪩�&�*!��}���������Si���g�*W���� ��l�5'��b��r�*�\(��yF�$�鴟4�=_v��=��`�뫕�����	Wk|�\���M�C�X�J,��'���>df�[��V-ۏYۏ���t�s�j95�_n��͚k�.7�@��h��R	���u텐�.�]#�(ה�^$m+x��G߄ް	����y�Q�G���2���Qn#�E&j��c�Ӈ��fx����Ө+���<j�o#��{%��]g�^gM�(��穭��ڄ.d�Y�b,��:f&�r����B{�O�6偘�s̍y�d�3����i�bN{����<1݃��� y���F@sWӱ�JZ���������ԥB8��uo:����ݽ�g�݈K�Oώ���|���+#L�d��PQ��R��17s�Y�_��<PrX�oʖ�}���V%�P]�y>������ؓRd�P��c?�1��x����貶����b�����OG���Ҕ5ȳ)�����^�[2	"�