XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������d������B����� yNi�m
 �3_�ml��5�P[�ȟ[�@)^i���ʩ�6���M3n&�&m�Ԥ����LE�c�Q�ʎ�a����}z�>l{7���b�!K��lrA��gF]����1����df-����/��^���¿Cxm^�r�T����"����`\�D���Mz��k�[�0˝���f�f���� 4l�B���<;�+.�Ɔ\u��m:i��lYC᠗��y2���d��U�s =[&�H�%���*�J��b
k�=V�j;(v�S
S�h������z�.�b���w@N;j��]��QR���zvq�瑅>�F
X4���Dշ��6��O��X�a��P����u�/U��3������s��ғ������K���hZ�2���p�\�Zk�->.�ᝏ8ʬ������[����	�5��=lA�p܅n=^h�
C���D#&r��d	ZK��}� '% �T�1wʾ�~l�ɖ���� �	&���1���B�L ֧����f����d�(@�BJ;�6\�����xlFV���5���W�k��E�=-q��F	��͔/v��[g��c|?���� Ʌ5�]� �z�\�sS�6/M���X��j���G'� 9e���,tKUG�u�ہ���F���V�txގ���0�6��X`�K<�Z�O:��o�ĸ���{��J��FU����F��F���o�5�0iC��ǠPB:��1Oj!�pG>ˁz`o�S@1��o�`�XlxVHYEB    10f5     490��ފ1qX�I@˝���E;�?W��eCk��R�B���F���{ �:?�'��5��k^F���͍�y%�q�׽l�����"�q��g%L�^Vc�s�m� g��P�#�]�{����[�����7���R�*)Gc��\r�}��$�i@�%td�а�]oۓN|	�y�k��TZ[�.�A�ѷ�K��}�Ʌkc�L�W�R�4��N��l3�Jq�܊P�#i�-�,`�x���L�\�(Y҂lK�gy���F�u�������zj$�a�y̸���v[������-Q+���_���\&��� �rŝ�8i�D�8���u�)*|��nT�@s-u�?[|.�̾*���1������0r�vO�>C��O��3����=f9X/�c�A{,��6yV�PN���+m��?�͓͉9ʤi$�R�йA1�g��hҩ��-L|�|����+{w�7c��a>�J5��]G}6�{�57TЃT�����:�C�W��h�m9K2�[�XQ�)	�t�s��^J���k���vsi�t���B���ZlR->L�xh&�B�'W��K��z;�Z�Qd+�ּ�tb�������]�nO�e8�e.O"v�㶍}��&�/��i�[>�vP;N�	e�A�����m���d7�ݾ��w=��O��ŋ�c���}�U��*���_��°Tz��M��(t���Vŗ�:�ƳQ���c]�c�1G�M�|[Rt�8[��M��WX���9N��N���D	2�Lf0	1�c.
Aں���p�Y���,X�+cQ���|v�!=�|��6�/%ůaƀ��]6��&���׋1p��qph����������)�0���i5ł}B,뷐�������%�x �L��)���M�
�Ԍ��s�|��I��ԥ��~.��Y�3+`M���=8���	r�TF�8hG�K��ى��8��˂|��Dd=i{�d�P�9p^�V�u`�����`�d��ҪEN��hT,��Ӽ��m�0�g�R�f�� ����l�y2#��י~�ӣ~D]���gӊ�Lֶ?�څ�RO�w���iK���(��Hǽ����tGl��9��z��<�;VS�W�&x�-4���=}�� ��o�}-���OC ���n(��B�#�]FS1�X�