XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��CV7�Cv�K� |�o����l&%`�^V;v~��<���?��Ge{ �#	b�D�<��A'uoƟ��Ԣ���v��O`��a~'��/JR�:~FA����hc?�3�J/��O��4����_��F�4�-6c���htk�/7o*�K)߯��?rf5��@���7u����j�����>����Dc,����|Z�7�'O�j�v��v{�E*;�N�����(�{9������?���嬷@F�T��'�yx��Yؤk�����H��$?Lb�;0f�o�ʟ�&�}����#j���t�d�eq�6���H��,U�8�X��Iq\CV��s	cL̀�����E��B"��G)�Z��+ܷ�v�����uϤ��� �$��B�~H�1��*�t��e�n��j&�VcR��d���rd����9^V�aݞϋֿ�^��qiy7di��i�Q��E��	�5�����s**mEp�؈ƪ�}�9�א� ��0�ʕ=޹�6 K�[(m��BiV���l�:>%$��ozx�S+x;��=/�Ơۋ}j�f��ܧv�K+G��۩� P�F�`��ڿF���]��	�j���߷+�sJ�I���ŖSZ��6M��H{
�l����iS�����%/�`kFw��1�?��` ��h����M�F�i�%��d�E��5tJ�ʊB �ܡc7��N.p�
.�]n��p�.�L�-;P���@]�²t� A��86+5�E���֢�h�C����-6���d���XlxVHYEB     99f     360\L��]��3�C�O��8��Y���F�Od������F�֙(�+�n1��S=�Ž�(����/��P��M4�4VO����|��D�q��pz��i.7�H�h�o��MA��G/^o0�v/Ef���?�Z}Tf_�>K,Ee���[��%�������"[#����IRu��-�f\�����[�4ʕt�?��V�k��uC;�e|>��lAS_Ց�Sk	*'�}a�3���YC+f���V���!��}5�j,s������pϬx1U«+a���4���/`C>�cP5H�Ƙ�1ݬ���=�?��^5b�4M?&�&���Z��
�G*xW�JbO�բ~��v<��:Jٯ]t��3��D~}}]�z���aP�z��z�z��\��p|�G�F><���]&x�7�$AL���ٝj"��`�r�I�Y���[�!��{��$#�����<]�w�I's�8���3�X�V��1�0ʒ����`֩l��&�ʵ�P���iPq��M�C�ಪ�3'mֹO^�J@l�;��Z[Q5���u�cp����bFY4�Eh3]�e.x����k�x���:v�>p,l�+��mBnJn��ok7��ELgP�;�� ]X�����yC.��J���~+��˯���s���¬Q#s��Ý�t��'mw��uK&ۍ�(x�{R?�P	2�gA��|��SK�Ny#a���)j�ڋm��T0�[��L:���߯_PE�T��ݷ�U*.0>���i����5�~j�ufvƙ��YB�3� X�HhHb���x�/���>�'�l�o��8�$��FW��@A�z�)O�U��}=�/(�����E�M�(��Fp�'&�I�,�