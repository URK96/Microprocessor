XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���=�H 
����B��o�F��@(iO����T�R�:Z��YYQ^�G-�p6H��+�j���^~n��ǵ��m�ʾ.R�>����D�2Ҵљ�˚�2dg�pT��N���pg����|v�OVREz�+\$��k���a^߲m~��A_��Ѯ���v���1@���L(h~�Q5��a���6�k�`���H$�sn>?�8*,�Ii5�"8�g����u�����C�O�dE�~a�2d���������w2.!�k;��4���ix�YxD�	��O����I5��ZW��)&��s2���q�'��Ej�u��6[��%�.f�*5��<�F��-�<�=����Zw4~�{��a[�Qq�)G�X!�o���7�������b�]��0���3 ��FY��k<�1}� ������y�<}8��`�����{�Z�F�/_��i�����x/�h���B�N�N ��ak�r����;Bʿ�k�:�õ���E�-�> ���n2A<"��D�R]��A4�a����z�;p
�&;jD��c^�ሦ>=���PEan���آJf�2[�m��޶�--����hs�bG��� C5k\#vIy��fӉ�<�$B4�;��� ��)�c�5��7�˴?�k�+�_�|�){u� >I��z�U1���)E�'
�f���ntH�x�?.@�+�YB&2K����I�N�[N�a����ڤ?
�e 9���G-�p��N.Jw���f1��?_t�X�[���XlxVHYEB     bbb     480|�*� ��ۗ�:�p.m:�Ȇ�=ہ0B㈛]QY%<�ͣ��C���2$����2�wF1V0��V���d`��R�ѝX�CF��$1�Ԏ���i�G���3M�D���(eF��݁$>�3��&����ǎR��h�ͫ^3�X���>���'{I����5��B��/]өtB}Ⱥ��ː��'���̳N#*`YV�N5Z�ad�y3�>������>�u`}H��+���	t
�ʋ��e�G����5�C����8���yG�1��^B��@n�K=ߩ�����Vg��ǝ���$eםz�x̜A@�wfn��ŏ^ۇ@��CHd~68���� �?��V�hP��:�5��A��l����8�FrT�=]̶�ݹ?!AK���6DrW#ث�D��U�COK���ف��uj�^�Z�4�l��CD7�6��~z����{�Ze���B0`����@���'7���͌`��V>��&��^��;�V�F�lin)�EG��I��F5�c`{�dɝbδ�9�9HL#��R�M���J��MWˎo(���dO1-q0
�	�ą�L|�����{�v�wC�X�,r��
0D��N@�jv�u&H�d�Z�v��K(��wx� �iV����m#2b�'��!x?���'=h���u���A��q��o0������Μ���}��'���ڔ�z��g���)s��I��̥'B�1X�Cj�H$����T���|;xD�)%F����O�;lk�����HB�hA��/�_��+�J�]�����c6`�S���y5��7}��=�z3/�v�u�7W=Qo��5��
�ը��D=��QJF_�e�Q����x\;�]����y����3��w=������E"���[^>��OhZ��S�������ƻ����jk)�;�=�'FJ7YFkѨ,2�&��XE*���Ub�`�+8��^h��Y<Z�9����2��
�p���?��B���B�(��RVE�q��v��pdV�^�I�=G�՗��(a�4Yk)�_��	?XO�p	�6"x�#���Y��O�׌4G�Z�i3��eT���%`�R�.R50��]
*��W�x9�#����o�1\S�5�H�5�,m��͊�޽N�>�������vB���