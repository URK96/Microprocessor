XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����A;T4���6�t�gBɎ�8]�D̈�Ā�υ�hp�>k�%+~g���8o?�^A���X~��u�����S�߰�!y�PwIg=���j2�ѱ��о���A)��W���'�c5(��W����U� ��V��c~5^wIN��lW�i[A��51ȫ3����ϋ�	q��<F)���0m���m���-Ϯ�W�y�?u��u7يz���u󇧭��5��ՀhJd��Zi%�PN�L8�3��LnoI}��IԪ��_!L������t�w-��g�Zz!M��Ǡ��<�7vccO��6�iو�{'����٨�9 )[S�`�I��)�	uˁ>�8hY��!p;��7/�B�-]�����3��3דd����9�A���x/hLR�]R�W�<�2H���#<��@�:��a�X���+�C\�4|�ф��2�n�S�.v�ǅ�%��i��wD��6'?��ᘆQI����AT��T�<�O�ߡ�/��c��ko�~�z����&zf,����H���'^U��o�n"��p����
�G�Nrױ�S�r��NKzE�`��&揗y�����Q �\
ۥ�s�����X��$�G�U��z��:���J��L��Ej��5{C��l��"μ��ſ-,ON@��k=���e���ì�uh8MmU&."���A�@'o�A�R�MĈ��ɟ�"E�2,U�h������Vm����T�e���������Auh6B:'e�h	v��@��G!�O��DV�+Qj�îXlxVHYEB    41a2     c20����w*�%C�?x��(N���h����8�#��d�z:R .Rc= 3�~m����%N�a����.�/b���T���7��������.��j�N7|.��{���n� �e�Jm�_�(����{8pu�,�eD�����b0~\��woI��c�(�8Mv�|a1�T(����	��릍��@�r��jM,� �������K�����Vݴ�>���F�{Cr��*'#GP8��H0��ul���o�#���젣a�M�O�*�\��y^�H=3���&d�ʒL�3��X��:)gyB�/\�&�rp�N�GCn�:u�tz,�c%�1s�g�*.�F���*[���\�C���*X��Y��RE���`cu��� ���t&�&D�/#��0��Vfb���䲻�V���檋����@n�;��q���Z�(s�M�$(�� �E��KZL�ǃ≠���������z�b����4�]���8u$k��.��_Fm؄��檜nD⩾�Tg2:� .�;F����uR�a�0�lRua�I1P\)f0Qz2`Tx�,�B$e�^� %�v��׻J��O}�����XA铱l��㛠k.���>�E�F0GhY4X���\H�S	hуƹf�����)�5�\��&Gh������V�#�TT�0V�y}�3
�VK���|�\��d��2V���SQ���ޚ�c��+����+��_߂TzC�H�o�.K�P��q�V��?j�/,V�.��OIܳ�,��t�(�t�dD�
��L� V��?+��;�8�1�̝I��ެ�h�n�׮��	b7Se�Fڊ+Z�����á�}��TF(�i�t4!��K�v�H�K$��E=�;����W�$zX�v��)`jE����E��Zϛ�M�,lY��-��[�3Þ�l��)h�=�BTXهh��F�J�j�����p�ۨ�{���'���n�1�dl�S<e��IZ7)�l[i���I5
(N���G���`�2r��}9{3�-�`�>���4��4��A��u*,�Qq�v?��pɧ��z�x��߫�x�~%�m�f��S��MQe�!��U�@��� ��� Q�5$b�T1��c?��5/�X�eW���������=,և�0r�^S�%l-!��#ӌ��E"c3I�K�2���I��w"�gh�?\�晋����Mv7�
��Z�XP�<�@MVJB0�����U��5B;r�FB�.��݊��P[Ɇ�b��hI	(�THi�ST�k3����h��A|�A8H1���j3Y��d��S�>oZ����8�4�	��a�1Y^g2��-VO�@.��;���)�ϏN���6�;aҫ���t���RtX�:���p#K5���J�iRhU�C�?�>f�ޥ�������a���΢d,,�N��+���Ea�U�c- �v�O��N��2zs�S��{Є��3���BH�ɵ��[�W�����&[���k� ��Ι3�G��!%�-�g����������������G�q+&����7���]�ڐj�.���S�2n� ���]k����L�I\�u��X�xu���Л�V`Z}���rc�޷ˬ_�������8��~�G���Q�R�����]*�]M�I�'�T�D�f�;�Z�xq��\-[bV>Y��O�p��dKi�L�V1ѢK�����x��/�N�K�JnO Ԓ �!�O���� �cmw������[�a�M[�p���m���	m���X��nոN�(W[6כ�|�
�
��ԛ�$lp�F����Dqr���e�cl��#)WQ#y��7*��d�׉�X��qv��$W����+�Id_�d@&��[)�:
��;�6�>\���`�L)�S$
���^�P�hM)8���y�Y�1���0��+S{һ��#�@�o�k�y��!Yh<��2��9HBN�z���_�pr�������6	�:wHGC����0-��g���h*� �Z�����ai��v����`y��f/"_M�ƅQ�����@A_�:5!�Cb��iz�(� �fR33H+�q�J��/�)ހ��`cS���F���x$q��hžLOL� bPD1����â8#4[��c�����7#�E�ʃ��㩸��q�)�s̬���d�>tϱL�W������B�qk�mm���M,4/��qk�n=�|ˊ�V`1++�dw|BM&g�h+pY���%͠�.��^eD��la���,-�u0#�LG�,��u��B�G�@$γ�i�q,�a ]�ؓ��L���<��̏.�[�qЉSL~��#��w�t�B�I��R�;[��x,�-iЖ�I�&��<i��9>��
���@r����V��ު�(��${;�z�6%z��p��B�	CM�ō��#�9
[_n�9%���9>��j�)�5q�xC��D���t�����*4�j6��2��)�U� �[8��!
��@������MQ��/�	q��#����<)\�QlO���&�c�XˬM��v��ʅ�J�4��7t�8w$14�����S��Y/핢��_�0�5_����yW~-c�J[��A:ir��$|��<�}������l�␨& \�s�'dQ`���b�Շ�C���q@�;c/B�-�z��44˹��p�� T,��lx��z6\����D#�wb�M6�$�8'�;h.��3��q�c�A�l&��W���>����?:Q{�^X�`˪�l=��jWO*%�Jnk#b��Z,�;���~H�����y�Z��$���}��TA���1�k��Chz�yy�ď*l(" 
�9�%8uM�4r�S��p��^Zz��xS��m[O{�r"M�����'mM��:��I��4��
�m�SDg(�Y��F�������*���r1j�ه�l�(C,�D�����,�v�(�7o� R6\�m��+�S�+l1�ܝ��Əz��Jr�)���'���U�y�I�K��r�`t8T�@��_�t�iǛjw+K�n���#0�����5�V��9^n�40v2q��\xy3�`�ǫ��������H&��P:C4��H5P wY