XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������s dWZܥ
�؁��G�1����y$Z��B%�O�dZ�?Z��-YH5�Wib����9�7ܩaƧ&TQ�_�<h@�;#��%��% {Շ*_�Yj�������b0���أަb�4A�'q揞�+{DLJ��o2E�Z������34�W=ږ.{�ЍM��My�����:�̘2(7�Tk����&�����!�	����ӧ2�Q5�8�3� ̶�me?�8B�R��*;|s��hy2淓�����.\��8<TɊ� zv��<�E������l�o���a>��R��@������9���t���䈻�l'z���2�@����V �p�q��`T$ZF�]���>HY�m��k����V���Y��S^���n1i}�X�Q��yi󰑝�-|��0��)7?˴��VK(�5i��Jq�FL	i��#C�׿�5d[ڕmŒ�%��0�5Û�Iy�������ڟ?JW��s�U�uV�}N����jRD�Vc���A^k^���Y=a��*��<n�*c�rbUX0�z�;>˘�>��f�Z��,1�*(V{[?d�fmu��6e�1�/�/���Q��i��_��QyS��u���.����/f�L�� �;nX�J�\.��¼z� kAP:g���(�D�cc��f����ӁC�R�qW�`S��e������Z"�92wf6�-��Ҭ�r�ﲒ�	 T9�܈~�)���M�8���cܿ���_�Iե��$������XlxVHYEB    2816     5e0t>�Q��m���NV�$��������{�)�Y�� �D
'�u@�_������C�{8��+om0O��,��/n�}G8r��ڷ�ϡO�?���v��h��z�������i��KC=i��-���*P��219g�Յ�yyq��R?���z.3!�I��7�hyu��X�x*�4Kl4�RصOI�9�W#��,��J-��Sr��*FA��>2�j��5U�N���MN
:(�A��J�i���]����L��ř��a��-$Y���թ�mP�Hk�Q��� �=��h�M:���\K�?���p���&j��
����O;�|�}x��X�o�K�����|J�j#n���p{���'a�~���������ٷ�K|�a�ү������J��Qx�,s	��py9n�~a���;:�� �X�*̄q���+�kK�LW�ق�i�yGoN,�H!��M=�ԑM�+����s-�/��o��kBO�J�K��iڎ�q�e������>�׻-O8�8�IɄw���ڒ�]��'͎�Æ�������U9`�jZ�e��A�Bl�1z�۱]�do[E�P��z�)�uG�O�}1=���h%Z� �f1S]L��xb��ݠhWō~��@�H����R �'��#� �BT�t�&��t�a����q�E��2\�q����'�s)��O⊢YQ}���ZtA�ljF��UĢ
 z��tKv0P���(S��4��2G�^-ŚzNnb��Y1�~�c��V������'*Z�F�,�~�
,ʋ����?�*�UנI��Ev����a[��4���J��KcY�����G�gP���rǻ�H��P(���~^W��Jy#��D�θ�p�ĭ(������b�0�u,R��«w�I��'�Z�)�^�����M��V#n٧r�vy��Y���f��Bj[��}�� ���H�E)���)dt��%a}���q"6��	4ת��Bo�P; �m0ƣ�5��#MH�jƈ4E��O2���i=PA���fW���c�B�Be�1������k�^�ɦ�0�j��Ƞ�|!kj�Q�zt�p��R�P+%�0�Nn�xv�رu�:b�պ)���/]3������w�awv��xę�).�]��8V��/���ʈ^��9�U;�Ӛ�O�p�|���vO�����Q�B�P�6��/@��@\v*����h5�Ș-c(��Wʋçxp���,����~��1�\E�c�l��z�Q��Š�F�=~G$��~���<�n���	��!,�n�0$5������VM�m8<����c�5T���*Y�%8J�.��� {:�Z���b5"+�NѶ *7sta�R��jbpk_��r{� ����4�}�%0���=��fC�)�H����˗ׂAV }�3�tvϥ?8J��� C/|g�Oc��y;kٹC�=���5d�9�i�z��T�L���K�^�0HTr�4