XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������V\�C�>Xي�Z�V�������۸�}�H������z;�s�74l܈}K�.:I���f�Tg!ƪrߋ@�֟Ov5��ޟp��mS��ތS�Ay~�%&�����!A�)E�q'zr����;�sߥ�3Q$G�+!j�T�Y�6�/�S�N�t�=v���Mp1`UY���lC4�����p���v�r�m�gY��4>���/�ŭ����4}�+~�����i���	z"b�$Ė- ��ɶ�m�D�/.�	&��<�6K�l>4W�&#)K���2��)�uq�?Zi�m�̤�������i�S�����.V�Unz�)�W-K�o�,�ԡX�0����[B;����5"�66�vL5M-������s�T)mN��l��#���-_��E ���Ka�] w/i��.���g`�
AKOў����&�4LU��jp�s6����g�XC8�5����fR(ǚ8�2\3�Sdu|aA���6��8 �L�vG^�Q1��2W� 0u8ҟg\Q�g��=
l%I��V
�|Z�.'~��F�Mz��0aX{��ry uMѵT��U�	���D-^A�[RE:��HBf�SO�e�D����%ݚ�Kܴ�k��Mc&s�Xp�&Ȃ{-�2�Ԡ>��39J;��!����7�-m\�B��<A�/�� l&�k��iN,I$$��m��C�]��*����)P_#b��6� +b/-lX (C�RS�l� "8FPB́}��`�/U���	�.�%	Pg�JXlxVHYEB    60e7     cd0_C���� f���}�e��lIߖa�`��{��|�Y^n}5�:۟?؊��M ��K!���T�8���g���eaֹ�ضj�`Xv�sd/ѐF��1�O��<i���d*�_8��e�s���g��y��G��&���~��V��dP��M�oY��d����t%.x)��|֮������3������E�ls�������F,��Goq�M��w{C���#�������j�.�:�	nԜ;W �;A?P�y!7�Z�:���"f����i�Ϊ�tRq�w��b�pH��&,�E7��^��s��ڸѽ�V`tZ���w�e	7�S�	w4�p���$�$��O����`MM��f\Nv�NPh�j�]��	�_�T�����xR�� i�-��ho��� d�j�PA���|����5`�]���t"�<��P�l�λ@�׊x�I~������F?��bs ]��l����
�O}ngJ
�u��9ɻlB��){>�i@��Ϧ�BY�G:����fA��a�,]�ȻK�ң�����,Ͻæ��DD޵��b�6|��������W<���.-��)��-�).ÙEɎ�<wp´2$$9��>n��*���!jqm �E�V6�����C���T�)�� G���d�q��t�$��ʫ���k�N�h��)���N�F�a
W�bV�w�b��!~�>Y����a�f���ţ՞ 8X�iY�A�&����;L� �y�8�Z �'��	:^������.��CQ�������^�.߀K�b2��C�hEro����q����"2X�[��.O,��Y����"��*>A��-���҄qHNJ��
'����1i���x�\}{c_'� 	iq���1�%������ds�Ř�d�M�f�=��Љ�#f�ة�t&���c��t�i�>Y,��-�C]|����o陡-��q������5�D$����ÁȞ-���m��'e���2��~w�РЬ���놝��qr�-U��H���Y. ��_(�� g܁s���6�4��0�����>'�5h]Y��+��ԗ�i�J�Wу�?zT��b�+{P~~K��{�g�s_�$����h����[�, �_�Fşl�a�d$��'����	[��x�����z�i��k�Նm�sĮ��M��Ki�f���������,����r�_K3\�,}�y��V��Aco2U&rl����*sC��-nuc�)j������27�w���W��ӑ��by���X�:Cg�Ŗ���l�	%cſy�u��w�H��?��]x���|:Ԃ��8�$T�!�8���+!�+p�)�IFZ�b<����\�6hm�����@6��n� 5�_^i�љ�ZX[|,�_&��g]7@�V��k���i�o>��}G���LA?.n88Q n����j��;�`8�N�79(������YI���a2�O듖�1��U���*�ڴ�M��d��Q)����~ԫKw����訏YC�Tv��W�*ȏvr�B�f vb���R�睢l��!���_sL�{�?h��<�o�1�ѯ�ʘ}�n�ʀ��=����|����~9�g'��6-s�i�)�k�u{M������ u*I���nXS�9I���n&�+�H�����')E��g#�s;0w���ux}�`���`���QW�� �h�_���m� �c�s0���QxH���<*�ٜ�?�lW�[6�8/!��w@��'����ƀ�� -����|��`�o���G[AD*��n~���V�2M2=f���zݣ<��
�E h��TX� ]ouxs���0�tL``�QI��5��4����*���q�CN���������y!%�xLՑ�hn�o[��hP��A� $M)�`知�0�ԋ�
S�G�p.8ՂC�Aw��Z�JN���SulaE\�u�zɊPa��}Zc�c��r&F��4�`llu����,�	[*�.eqU��R�[�wO��OgN �
�w�0%.PDA	�n�0���x9ԙb���$����n��+���F�A��:q.@�ӈD�E*(���(4.ާ�����g��5t �Z��Hb���س9�l�?�v�BlԮ8�� ��'�_hN��c ��O04w��Er����T������H����D�6�ٸIВu���4���Hԕ�|��Y�=�x��1H$41�GS�/8i?߫8�b����`��\MlM�+_\D�9|}��ټ5��Cy���aٻ��L풞u�<D��5�${���$M����
�����m 9�_u&�H'(�li��Dб����]j�P�)n�b�?!]�Z���|���y&�����A����K�ڐ�c�%zB��}�2C:dB�Ŕ�r��ͅ�6�FU
��<4B�2c@8�&���\����S��������_F֔���GA���
� ���DTa1W�({��3�K-QXN��d��B���S�U���#4������xv펫[}����Y���F��{�;N�$��r�<u����{�K$ ��}lj�/�돝��mU�t�nmTVR�3�J\�j@�^� h��6�R����K�
&������4���\0�q�W,C	�A�W���B��"pn�[��yճ�T��b[�]���Og	gǐ�뛀��ݘa�L2�9��b�	��i}��u�g����9��:�f�x���t
�����u�d~gC^��IE\���9�;K��tD�p׽�'z#ֹHE�c�q9 ���*-�rU>D7*�� 
�����0���pL?P���뫔@$I�b&&9H6A�f�,F�{$ @��N�j����3��v�r�FnoA���:�[��TrF����Μ��j E���?�յ�2쾖��E�R*�W��O��s�W+SƯڤ?B�����drO�Ai�s�d=ŕQ/�8���̞l�k9QL�z42���<A�7���2�W{6����0X�`,N橵G8Fb7D�̺B�Q>�ʵ)'��-�W�E�<������ig �@���(��\W�$���I���qwf�T�C�����ӣJ�-�v�l�G�?Ih*w�ҝ�U��Y����8��`�U*�I����*^�(V���e6�*����0��Π����*u���p7Ƹ#��˛ň������Y�i��?���WΖ�Q̵��7 +z��ʙ#a����u�(�{+���FO0��(