XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#�0;����u�\)��?x����������M�L:S⤸�Q�-�2�V0�1�����Z��)�/��e՝
��ō�k��R\YTA���(WG��8VV$e82D��ƕ���eY��Mikw dl���!n��V����+��^�jo��4,j��3�8�B�]C9��Q㚊��b'l�3yCf]�:��W؝z��L�ٰ����[#���zk�W�W(�9|̶�Be��R���{��J6�;6 �i��Y�gе}q�H�[�R��[��3�s�n�E/�H+���e�K�)�ri�B��	��`a$�	�0i�oy���������Xّ��
/�,	������(O7W���p��Ģ M:&PX�Vv�D�.Z8���~�C��FXR���37���{�7�{�F��r���E\��;�z֛�5�ɿ�h�@�h>`MQVp`Kj���ݕ�Y��NH���i�tʟ0�rkҔQҙ6���0ٶƍ���Δ��/���+B��z5�?S�F��U�L��?��]��k�dM9d�����
�Ysܺ��S��,B����Ū	4]�\K5�0��	� ���Y\]�f2wZ	T�n�F~�"OF'~�N�y&` 
yj60�M��
��H�Z7!�B��C�i��FLAd��h�V���l$#�G���fIB�B�]T��떭U��ӧ%�S%;-�׬��7]}�[@��i4)��R����W\�:L@����T��i�F� ����M�����E���DQs��}
,#��b�T��(��=mXlxVHYEB    7945     7a0 *�lRQ
�'�\{�:.�%������6�R�z-$=�Vu�ɔC��Bk��-a{wp�3pѤ���2:�k�ż�\eP����M�T�S1FU�p����'�xG:K\���l4�<{5�r�Ä=�<L��]��!H#�ޠ���R�������[�����Ȅ�����~>�C�%Ju2��E��*ҧ�Kd|cm�b��T������h<�b�E�f�V��*��K�m��b�.�`��+�o��)�f�5����e=�+�g�u��#?���K��fŜ����vIZ��Aܾ3l<҅p.|U&&��3�b@s`z�:�F������e�%g_�B�Q�F7CXp������>,1�CɏX��yW�6|ۖ��k���a9\��b�e.���Cc�����q���ᢘK��%g�^ ��9/?ӅLEq`sU�G�MbG+C����4����O.�oä����Ao��ncRچ'�E���$s[�_�)�y)�5�:zi�{�F 5�@\�qwA�Z������:��en4G*�at/�z��Q� M�q��ۃ&O�VD��kJ�a���s"{���6d��a(�X�Ȗr�t�W�7���^Ze����O$V.oPi:���2ڛ��MNS��F��#�
�n:�GN�PQ�&4(�.H�A�X�Ju{.����2r\�[�񜹾�W���s������9�#z��n|$>Qm����Wh_�Tn�h�G�$��9��_7"����{�Ӟ���m��/��kwy�QɁz�����/:�(wXx�7GD�I�e��إ���ѭ���v���������!�E��ǹ�6��=�j�� �=�ā�[�m�烆V��n�
�F����7n(��L���N�q�r����0�%pMU�HX�gl�Bo�8��Z�+�#���N5Z��r�����Ŋ��db�e��X�C�34���OZ\���'�v��X�~sc�zՠ·���g4�.Լy8D�WRn()3cp�}�@d4&c��~�Q3G���W�UV�����٤���k3�@:�����Q���[�H#S��Y`f�f�\#�O�np�����k}�]�dE7�j��6c��p������f�sS�+�'��t��U�����=>l�FiE����+_략0�A���X&0��m����G�iM
̻�tJ`jb�<"�F߮c�v���lk��	)Y��L`b>T�i�(���u���\�bi�_<�'�AH�[�^�(�x� B��������6o�8�jn�~��
G�/a�=J���毨����W;�V���@n�%�q0"�� &�n��b�p&x)U��X"����A�
�hu�]���QM��$�0Nw�	�3���5E�C�L,6b��4=�i�r�\�1=������,W�5��p���=�pr���F��5�ϲ�"	�x_9��Y�#������s����gU����qS�VT��z/(����ʹPBw ���dP�a��ک�-t��"��KuF=�Db~���2��֘�OS]S��sN��Ò�Ί��hdG?�)�2�N�3��"�_��Ō,u2�����k���7o,U"�|��ڦS'������9��J�Vxݗ�Bknb��S�UG�pj����0�"v�.0���-�F�<>d�ڮ��4��E3ۀ\l�ܫ�~E�2��Ds�%>�:�{��1��ߓ?ȅ�{p��|oqS�Wk��P�����8`
wȣ��:��ėy\�QcA�үlT�%�a��3ڹ����>�B�z��%~�o�a"Z�Å�'���!<�cyO-N�-R"a�N�#����T�����U�����W)Kh�4|7��}}EU��}��ɲ����N4�c7��u�%����.����=!�y|����.p�&䗯zn��;)�a��)H