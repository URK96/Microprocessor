XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��s~��� ��FC��?2I�f�w�l���bg�-L=٤�O9@�c&X%�ݻ��s*�������R��#�,Hд�̱�T�죹�+OL|�Q(�'�0�gT�TOb��@�~W��2p�`�"�O�̦�D�`�+�����Q�B�`�ߨ�1T�߈6|Ie9z����/��D,j��~di��$�}�ᶇ蕸�u'�j���h�<�*���U�c]{����Oy+���U	�4e3-D�EL�F�Mᢛ���`������]����fMW7�ȭt`"��^��ʉ��ڎ�h�!�BMŐĈ��!z�6O�)��0��G��<��Bt���#��^�n~��Ɂ�ϊ�M�,�o�	�n��&��c�#?�x	�k'}A�i ��I��ҹ���%���������fI �@9�5!��{�Of�2��6`��YJ;7�rF���Q�ɟ�(�H��[��U;�m���P�,���i4��p-oa^�TYj��}��}k�_���=�'P����o��n�����wι( �5�+��7F��IIk�T`_����ՎJ��{I�8^������d��Uz(�%)}ER�� ^�.�=���V��E��E��Csd�_��%�*>�b�/��ۣ;c��Z�_�A�Gۼ�`1
�\�l���*F]H���1k��\(������l�k��5��D}�I��G�>�~Jn���$�{+����U�g�1�݅u�G,W�lel�@Ok&x��%
��� ��M|9���9$فڱ��t,� XlxVHYEB     7d5     300M�Ƈ���|�E���L���RTV���0�Ȓ^��1�Ԥ�dB����l�~{�dy�bxj�_��H�{�w�c�l�! $J�����g�w�e���K1a�����.|J	�s�̆e�b�ͳm9�Ϫ���y~�,M��$v�����o��-Ƿ7�S�A�f�~���wDA��_�����U�t������+l0�(�2F�|z��D�.b%K��F�2Ȇ�R~���w+�;s�}P?X�p�[@#�{4K�e��Q3��
��cn%$����C�h�diaV�L�t���e��8y*A��c�'���X�wI��_�U���8����,���\U�O�#�	M��:�����n�^����sV*¾z#�|?B�74�2���Wx�;3���*�Cǔ�3�껵c�M'v9#��T�]yU$;�^lpU�D�vGϦ�4�A
?��zϽ����.D�ǋ�c��L�4�?�m��=�DH�6������A���Gv��_]{��9(�}�U�0��s}��j
��b��wAf��X�Z�>�!fi��Y���Ƒ`�(�H�/N���MN���/i�4o��e�͎rM벦�� ��i-���Mi{�K{��^������d:��n;��~�<�������!ۘ3c�~1���T�"���Ü��A떾���}x�������Jf՞��;�4�ص�$�M�� K�e�!�1"|Vߝ�$;�8feY pI[���j���$��<)J�#�`�0eK�T��+�{ӗ� >��