XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9\��1�3�l�@T���ϴr�,}Xδ �WS9r`b��JGg�9�FE�e>�I��mJa����_��)��ˆ�:�UQ��K9���y��ۖħ��r�6~�w��=������ڔ�OQ�}k�@?�>7g�F#0>I�j�~L�t���_YN�ڜ�vq+�ی�g	8�*K�°�Ws۔���a\�M����ReC�e���ճ�ծ�m��^����g�W'<��ɝ���{��މy�����n�+N=�#i�9��H�r�M�,�u<��>�~�3���g��-�����N�#�I�D��ɳv"��rt����{�Yϴ��~��Q����Ql��s�T�/���~
�r�d=����j�e:����\�pm���v�H�{e�΀����%#�|Q����@U�s~�C�z4�eh@S8�~`����q����1�Jc�n3�pU��ev��!�KK�*G<��D{����N�Yj��뙏��y�aWm,4�xf>�S�c��U�e1��Ϯ &���\RR�쬅�}��W�[��@�,w;ϒ|����&C��w%�˸�z����*g8�ȫ8�M��2���g�:����kC�|����B�KI��d�9��O`w%��`��~�C�S�mA:͜�h� �E-q�~7�K0�+u�X��T�����6��D�x�uI�Z$�"~����Xh���0+��:� ��G@R�؆�E��Z��}��6b��j�n4,#C�.	��k�cq.J� �\e�ZB������9�j�XlxVHYEB    6df0     b60Vi�⸋�8������ER#h�g]�'E���˲��1�
S��]/F�\T؜5�<�q�^ -�Q���<s�q�,����ܻ݅���?�Z9FpJ��\��и�	u�����P����g����l��{����1��Ip���N�����%���>�ccu��i���e�X�F��9�I�Ҷ0�T�į�Tц�V�>��=�̹��]˂8��ƬV�eJ-MN �3r�"
�R�Y���^3r��O�����Vu��`V� W1t�4 �P-֏��H��Ml�·|V����.	�ZO��i�p�e���퉖O:LF�X�ܬ�~�����m��tGD����C��������)�k
)�>H宇V�l%%��4��r�}����}�1��,��o�
tR�k��n	L߱+�rR���X�'Ǵۍ��G A�6M��3 �b��&^�5#�= �~co�S���)����r������;���m{p�)��4r5e���A�/�c$~��,��2Df�����D?��s�=��n��D�t7�����D��a�L�q���O�����%���s��!�Q��\�6��q5N�PT˟�3�4�<��L]GI�E�"~G��`�g
�����;�N(0׿���N�қ��siϺ
��r~�l�~0�{��H�\#�7~���^�2�"$nilɘ�7�#SN~(��i_P�7�R4�}��s:ɿd��R�A��&<9���hűF����Cmy��C�gѡڠ���bo�E�ӊ�"���<Q�#��lo�yq���@��'f?w��Z����l�R��쨁�]a>�(�@[a��D��Q��o��!0��q3�p�iUZ����Vi���W<��nG�X*���J�R��2~�F^����@�I�i�Y�?��sFC�P�[^Ņ��s�풌Q`���B����'@��c�H�P ���w}��Nc����yFh�O�}��^����3�C)J��oQ��@sc��/�I4�<��A��,o�߱��0(SN�_���:���'o��^�)�PWe
�F���.�$U�����G�@��n�۵��*���f��[r�۵�)�/�|5�݂�P�.����R�#�T<�IU�pD�Zq%[�4��P�ft�t/��ah#q~WJ,;�8���T'��ǀ0�*� O}��ScU�쯻�<ۀ�Ǖ?y|�e^@sʋ��+�)����($w��f$0������$]��+�@��6X+`\B.��
j�#B3� ������HJ��i�L+�lu��!xY��w��k��Ԣp4�B��h�K������:����Hj��j��%��j�6���\�m{��L���~뿪��D�Q��[�9� ���1En���f��)3��^�#�('sq�6v4��IF
D��`>CP�}+�<K=�Nm/��y�cI�|��Q��w�[��+���c�NEn�������̢�ad�BնjO<`8Q��T7�W� B��b��םm9����)�.����l���k�"�I�/��m$��H0NO)HA�G9�3h���@f���R�{���-��F' Y��\�Gs���>��2�4�����������J-���hl��ۤxa~v�[*����kstW�����w�:���`i�Bj0a���#F��-�H�w�iN٨4���hj��`$�K�A�Xb�3�R��g��U�ɻ�*Z9����-�}�m��X��x��G-i|�����3|&��G�7�0���OV^eO����pt7�n��k5p�z%�k\�b�YŕD$�.�ݻ��t�B:q���	���NT�@e�݇��sԳ,�F!�u�w�������_dq7_���1�=�WCc/��Hԏh���FG��T�ޖ���%T˪�}�0�R�;x܄����i%�`���#�RZ��z����~׵��݉J�F�O(��$Z�*��͹��CVD��{��,o���ܬ<S���M��dU�nw��A��%!��7�<䍈wxW�L|�:���F_V� �kM�+ې���OR�p+[��iO�� �4MH��W9B�`Kq;�Cdͳ�,jI���=�L�+�K�֎�K'���S���(h�3R�8�V]10��md�����-2��-��Q]·R.[��2e�ދc�5�W�+r�gh#���f[�5@t�78����{�>[<}Ȣ��pk�P���i� \%.�['vt�2�N��c<�)�xg�ăI+\r�����L��\Cv�mh�1��M��ڻ`���k��:OIZ˽fy
�	��0�Չɑ������Y�GN���n[>�,̈́!S=Ȗ�|&�u�6�eɸ^�?���B�t��5�1��<l�����?�ED8:!Ӈ��Q }[�����7vKS*��T�P�t�',\>��e=S\0����$*_8��M��}ݓo���t��ʨO������g�7���г���gk���'����d20��:�3��p�?���6a�+<�'cRL��*^>X"0�2%yZ�l�����i9[uJ2hb�\�]��d���Y�Sq���2)[j6�@C�ꮅ:�6�EY��(�����5���$e�������!�Co��xȘ4U�Ƣa|v��A١n`��ɤ�L�T�+�rH���k�-o����ER��Drb�_0A�:Q��q��$���֝��x�6�݈�RƤ����tJ-BcE,��Ő����xl�_�z�o,��e���Ū�9�r�)��P N�OUm&[��9�2l�
޳��o�:���.�V�Ø����T�р��=�Q�������4�Ƽ-~䑦�8�����)@�U,s?��Q\	����n�f���>� ��m[ۯۨ�