XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#y�*(GJ@I���������0��+3�ӇQG�s(b�T�4~tT���GuP��(�k[g�x��f]�[�u.�@A�	Se��gx�i̝�sss�Վ��#Ք!���x'�i|(�d'��(V��馷*����n�/�ې���n&�7\�q&!b;~i���.`��Y�)4��L?7�����N���=T�����\�A��u�e��H���j�"/���Ӈ[�L��BC�n��U�O�F�X�w��S�4m�r�?�_����13tShh /RHm6T"����!�n��_��6Zn�xlÑsܫ��(�n��u�f>��9�T@!v)�	j�Tc�&̺����םz�5�	�@ĕZ��t��7�f�l�Jn��*Dn�A8�X��V�F��	�m��ʣEOr�����v�OT��
 ��h�6v&���B�ި*.��z�B\Tq�f�4�y{g>�+S��E�������O!Y�p�brG3q�T�ҥ�b�w�	�F��H���_R�˨3���4уƙh��g�>�d�i7��=#�'���������&�Q!4�T=�K�v݅�s�e:0�`&wȂl}��䜰/���F9�>�R�w:�Yig=�ۈ� �������?��Y�0*u�*�nc����{�7����>¼W]2?��(b]��i��D��d���H�9!�@��Lh&�0!`�W�v���Y� �܋r(̴�X�4,���� �4�`�M(aٜ���!��ҥP%u	�"�.T8Գ��5:w�XlxVHYEB    3541     ca0F
x�_�<���X��_��ݒ޿\��ZWv��& N�l��,>��;	��s����G��k黵�X���5��m���ǋ��#����������a��V�+�����s E�|)JF�v�Rk,#�+�-�z��@��u ��8��7�kӔ�u�3 ��ܮp���������o��7Qn���s�� J���^b >P�q���t :v��^]�@���j|������^�ܥ��������RL.��
�;f��@��X�I��J�א>_n�U^u�ы���;�Mfō�uځ���mB�惓����Jw_����NG��5w�-m��D����0]܊�!��k��'tQ��ш�\��/�?�e���|�Y�P�C%9K݄�@"�Y�]U-J �0T�
���d�&�Zec%\�dlR,�磒����q�	B�!P[$K��k�¡*��2�O� ����ƅ'"��{Ėg���cL��~��+8�M�:\.@ܰ����u�7�-��-[Έ����O�ߡ�~r5?q�W�>���������.�P��#� #|!�'�Q9ܼ+=	u�n����1�7��v���n�CO���X�6�;���@��mڠ�l�|�9���J,���S��ҔR	Qo�7aY� ��d����G�����5t �zW��X��[%e��M��k$ ��N?�~�7�����E���M�T�d'�f-��e�A�	L�Vl���x-��8�h;M#G�u8AE�D4>��Թ�,�Ԇ����Xnw<����%�V��ޭ�I��O�To	}��N�%b:�D2��8�QǤ;�<�f��l5�/��3xD�u���t�&��Y�@�-��IM4��֡�_�U s���Uw�j�� *t���v�&O�	.�����􂆃����*�x��`Y��H��v�aW�h���z)�����8İ ����)����<��9Z��;i1�|
����{L���ʹOx�=�k��S��[��Q�j�����`v���E����GW0��P:
e�Ɣ��;CwG�����־���蛟H�9@�sXw��źF�}l#����Y����n�8-�F�Y�`��@f"S�,�-TL�B9�F�E��Kmd�8��|�b�<q���WW��c�*ۙK`�?0���ǘ��j|M�����*��a �`��c8L�L���N��-W{U�����Nw���̫�]�$���W%�c�������7^}���r�HՇ�ϥ��`��FU��<��D�/� M����ɁuՈv�M.=���&�q�+�e�V{���:�iY�t�
��t6!�;�MCe[Vį8 �6Y�/a��eȃ3��EmDW�k��SA=��8S�y͆/`���3���:}h�f���j����t�.���0��> ZX����0h]�V:��Sc��s��/0��n��,Y˙/�V����L� ����Vu�9�2�Aa�c�1��l��4,�$z ��I[Y{�	Z[�ۉ �b�Sux`KR�ͰB�OKâwK�a&\�Rudbx`���nÃ��јi�+ƿr�n[�NI�����(��4����5���Y
�4nڤA��F��m1R!���P�L��c��v~(EQT�6)&X���?D� 76=j �^�jr�l^$:H�	?>V!u��e�ۙr�n`�q���w�W
<��?���n����:�|��"^�[����7����U6�^�k0K���kW呄B+%�t�v��~�|��ӓ�v�Ɏ|
E����9(�`߁�����{�]ܻD)a���� %ݧ�-�$�y����Ǜ>@�j��1�$n�)�,6U<�_YBh�_��4���'��^�NE��z)x>���yN�"1G��XGIR����d�Ǎ�-�7(o$lšQ[�s�c��D�yH�������N���3waBU`���6F-����=в��aS�kM�����k=�1��T��*��K�)��3���VX1�0��"9�/qy�_�I;-�k������>��gD�%����X�� V�e�8ŢnQc�&����`�� Tyu�1�q~���v
��'8�l��?Y�t�yu;�	���8�Tg�Ù�r_�xgvZ8M�IkN;a�H�^#�6Ě��ei'��T�'V޾1
�Ͼ��{#��a u�Z�2F�+N���k�c�c

r��5]!8���H.#S
��=U�M�{nywD�Or����u�ܻ���Ok�y7�v��2�7�{���I�^�d#�����RaL(����y�Z1cx	3�(�3vɑ��Ƹ��N
I���m�����[X���IJ�!�:��@��V��<DHK뉷U�.Vi1���Ń;�@��ձ��M��.XN���3�D�'"F����e	�P�8ƈ� ����p��Ih#C0{��I�󋫸�o�
m|%��T���7��J/���7a���l�Yg�w%7�(dkN�Mt#7��F�8V��� �}�Yb��CmqN(2�Z����p=r�A��駂7ʬ�2��7���������ս�O��� !OX�;�~<l�8��ʌ�:����|�1T{��{��GTHðe&VsqJ�F�S�{��D+�ǲ��s�yU�Vf�c�����\��
s:I6Qr=K�b��z�0�i��zD'(�m��Ot Q������O�ʷ�F�2�t��u���������A�S�+L�>�y&14�K��-S�扐Ke�&�T�$:Ǒ�Y=�2%3�ϰ#H\'��� �Hj������xq���ow���o�X �[B�d��D����7"��Z��b���۩��ӝA���6{�D�6	�&�����,��k&E�3I�P�>���h��Q�|�S�[���S�~p�?���E�/7������#6�h�i�k�t�	f̺�&��q�<n���X�����u��@��[1W�*	=����^���ݻ<0p���'��W�� ���`��י����8�,tܙʏ�6|qO������2���o0���\y�E�,2:Ȟ+1gd��Qp���*-#e���͚kbEl����g���U�0�tgqƴ��Ç����#��b9�UILcN��|�Z!�vc/�6T�7{��MW$����u�o&�ҏL�41�����X4s?�Li�np!�j�M��Cr� 