XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<*�)�'��и^&�{0u��-6�Y��9zd/�n��!dr8'�]\��@���"���]W�u)�N��/0���Mi)I�X����6�|���,�iX��ԋ~-�by��g��Av|�n7��=]\#�q>c+�
�z�#���X�Ϊ�M;77�Pq�3�w�����gbw"�:���T+t�Mѳ9������������9���=��im�>�� �������Vm)���a�խ��n!�C�ѻO��������0C'�$���>}�'D������8���ʶwT��dS2�\�e?�xd�����QrC�{�Q�l�J"��'��Z��3��.���¤�'�D�W7���1Z�pc��-6�1���e���YT�!����4mS�q�$��`͂��լwސ�ĲU��a�uґuk1�+����/�l�������H��y�?�N�Ů�8�3�c��#�ʰ��Nq�6"e?la��cB;}V���,M �b��?�·�������]�0%a����ai�	����S�TZ��j��L�F��1�-��O
[��Vs@H��.>wSz8�6"��=R�/�mX@6u9m��%�ķ�3q�$#C�l�'NJ���ʀ`G�|{VW��a}=J ��I��}d�;�q�s6DЕ:�K��xf�2s��q�/��jg%A�1F�b�c��<@��Ƌ� :+o��h��n����?��T��bW�dI�'$zx�
�.���0?�Q���c%ng��b������`�SXlxVHYEB    9944     fd0�vۛ8���b���=\v�(>˷� o�s�A�KE[�!�� �R
��]�ė���+A@8�0ƥ+%hV�G�W��A�W��2$��P��e�����;RU[.q�q�}2h1�W����ʶ�rD:%{Vٜ��5���e[W�򺴂�cHY��]Y��O[[�^�
v�&�
���ǂQ ���X��gq|���A b�Ѩ�����K��,7�5%Q
p������<��A	�̓����8F�h\�t�x�_{Kedk�i{:�����C�~JvP4xZnu u��E�Z�0���	�lYd�>�c���G*&�1<�vkZ"c5ܺ��Z��%���%�3�1V��%�_ի�g�\[&=�O��#^N�G�� ��^L� ���3~�5Kx��0F�>yz�>�*'������r>׿��ƺ7@��l�)��ez��2OV ́b*Z��?!�N�����#e#Uu(��)���<�M�N����g��+@���|���[E��1�|b���4�.�q��H��Q��m��e*���Ay�˕g��Ӟ�_���bsj����=j�|X:䬞6���B�ܤ\ -�ݢB�HUb����r�ݸ%�G���!�"2$%���m8���\ۛ�u�.�=��(�c�4���g���BJ���ipܼ�7
;~F���88�/�ʄ�:�}����!�t��;ۊ>���!�h���%���P;�&���ܭ�$�a3R��'���O�TOͯr�(���w΃T�krh�S��B�)3�*� ;���P���Q��c�.����z�&����
�e��(h���T��mg�H��wٔ蟩�aq�����&ݳ�h����~_�3#�Q��YΖ:���k��<�W�����`5��.dV9'�?L�T�~u�8�w7E�_��C(��� ��V��X|��+}!�/�y���C2��ͪ�3���ʋ2����5�~u���4�]gp:*�����喖����Mk&O�.�^�}@��p������f��U�k
Ϫ�n<�+�n]�p�.'�������QPA�͛�2��۟���/ǀ������6�* �	��=^u4�m�.ޓ��Z,�b_��o�T�$*�V1�A�d n�^OGp�R�H��O��k_rs�N����b�-�&�*-d���3�@"#��c"R��?)`�le0�]�P�5B����;��QU/��K���U��r�ߵ��¹bCdΙԓ��w�meW��\��&R1�uk'ʪ�XB,5���IʇF㾱��2���3@��h��~n=���Fb��ʮ�	��������W\-��8Ҭ)J�ub�UI��@Lx	.S=�z���]N߸��a��Y�ްL��o.��N$덬���0���g��R��WB4��D���K|"�4�>}n�BZ`k�T��r�-�|�Kw�n����P���� f6Р��fچ8��A��[dv$T�osf$@녎X�ri[	����UW<uQ���:�E���R�^�M���Z�P�yG�*6��7���R�J�M4�~�$y�y/J�%���r��n����O�A���ʬ0�̨��@�Lբ�s��݌� w,L�w��z�L���({�\ՠ6�l��quEȃؠ�P�3�^�p}(�xȪ��쓝<ԛ���DE��醨����`�R,�8��!�����g]9bX��}{��'4�i�A�����8��Z[XU������!s (��|]G��Ƙ�wb�'��9+3[dO�{�DX����S}���	�]���S�·�i��
��J#���0-�0�-��6��s���O�0sm�j.Mן����e���y�H/b�k����:z�L��_;禮Z��e��Jd�U�Լˉ�2y���\0�$��T!��":Ts�G��y��!�1�����:Ӕ��'2�G2l��)Df
�p��/�S�v��-:�����z�q��l ǗrA�2���ȕ�2�P��,�3�EI���P2첲��RPoEw���aŢ&������fb
�����v�ǂ8��%����ԅ�����F�<O���2�Mx�mE���˩�2��uƎ`^p��7B۸K��1W�Ӄ����P���Z:LF���@�ة�+`��:�%uuQS��k^�),ƿ`��,��m��t��R���b�!���3sU���U�D1Q����b��b3�j��H��s+-.��5e�G��!��>�)Z-wӛ�=�p�nf��h��Sn��X�1�A����X�r�Jb��o1���w���<�.��ZR��I�S�0rn|A�Y/�7!�����2���Um� /'x\D�+�gE{��@�p㍾�o�ZӇ2eʚr���:Ӹ���(��5��z�/V��\V��m���`�OhH�U��׊"��ۗ�%�܅��E��!ѧ�O��Q���Rt�?�u����xR#Um�w"4oi;TA�,���8t��Dj��H=��oީW�
����ֳ�Z������O�����
���pה�;OL.�.v.��3>�V>� "��M���/�(�����&��N+l�n�Q��Ó�	�}Q~�:���Q@G�$V�ߘ��dQj�:7���^�(i6>�	V�,�9H�EjN���@�ǥ���S��HY�é)��2��OK'���m���yC. e>����2�$������@*@�m-|��NK��(�`Mqu�g��#���a�*���v$8�(:��Pr�*{5's"�z�)u{e�`�=��h
���n� n���R �k(�3l˳F�z�G�.�^�g���G(N�~�V莵��J�m�1j^^��'ɠ6��.:����y�#{�2�z�Ӧ�Hվ�Zf����Gi`T[��(�bog�^T���Ivw)>�_7c����$N܄A砫�'Yɕb^�?�[no�n�@��� �G.��?K���"��}�.�m��7�b�)*�B0�Jy�`T�\yᩮ� h`���"�qG��jr����'\�>rA<(� �ƻ�g���F5�؆E�F�w�6�Z����$�&�ԙ�BƾId�I�K�t�3���?�p�z3�"���l�P�r���ӡi>�xI.�%m݁'+�Q�8u��\[QT	�
�\�؂�$���\�X�ۘ��'н� �X�-����I�,:��8i�;L�4Yr�ژ��>�M�)Y����xR�2nw��)QF`���'� ���{�]�?�Ж��B���йb��z��Z�t81'1QZ�z~=ʚ���񰳠���'�
I��A�c���i5�_�4�d�<�ޣ*�k��n�D�ݽ�DC�ΧuS��H����(A�g͸���-����<[mMY�zۂ���L�i��o��Z�/�$��bJ��T4�	�N�ٞ���=�p��
��_&�媼.�a��K���M@����v.�[�Q�aZ�!��vߩy���~��k��fӕ�����P:�(�K��g~�$�ղG�7Ub%5�`RD�ǎ�7W��Y�����>��5��R�O �8t�m[�c�46�q@�v3:+9��'4��w�4��ӓyߢ��]PQ���M��OF<������ !�Xj��>O��Z���e1[ �Ƶ!��Ų��7u+L0s�O��B�ˊ�(���&�f�ꐃm`����ϡ�>P����t��}��n�%��w�0"Ѻ{��`��rS�٤I7Y�)��&9B$.XM�B����
�?Bb$�ϊ������F	ٴD¿$k|����ub�YtD:D�������Mm(���Em�L�6 h��`��%@rƋ1MjƢBPg�k���zn�[�D�1@�{�)��^���S��&ܛ&��Oӑ^z�����(�Bt��DI���9Ϧ=Q脁����K.���î���oUp�L�Z�mNuqSs��vh���>�=ćC2@m��t#=E$o��z.ڨQ|D�r��a�МO�ǳ�d&�'��~�k�<:��=�	�z�8���l�駺���