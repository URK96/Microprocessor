XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E���K��*G��NLس\����_6\l�k��J��]ԥ�h:�j0����x;��c���i�St_�[fk ���}��KIU"[���k��%0pN&Ǩr�m��h�e��xW�uh?:M�O���������ճ@ԠbI����v��o��_-����z�!�J� d�e?7���P²Md��xb����Ma6����>�������j~��I��-�d���4Xz�D?�Řv�!g��)~�ak �~KԿ>��G����-�f��l�)3�T�璣����4ʼq9��l��Z�� ����;w�^ �#T'jK9Abs����E^N�����c��E����F���\� ��v�a0��e��z�]Wƽe-࿝��((����2��S�Z�a��s���q���'3�,36:�ɜ���|��}�,��כ�xI��-�ȇ�Ta���}�����<}ϠE�"�������`�I	Ȁ}��;����Z�WEm�^l|#HR6<s�Y�	WY��|e*�^/�ף 9�&��_�"_/Z��W�ñ���B6�`嫺83�\��:��� ��'|X+8�1s�֞+qa�n��o,u�`�/�,.�U��E�*�K��>5c~�F�l��z3�8z�R?�y�����ksEǹM[F��9]6#���I�̥��!ţ�T�n���{�~_b��!]��FnEo���{�DFVBcc_��\�"�_��xYǖ^�٢?���$Q�ȹן^�w���EB{XlxVHYEB    3a15     d40݂o�K{Ɉ��o<C�b��������f������Z�su���ې\�F�6��Pa�?�H:��X��K;2�Q��V�#��C0~k"!N߬��"o���2g
]gj��Zz֕Ì��t���p�����뒢��w�ztH�.N�n�A��l�o|l��Htɡ�:�Go�H�����ɿp��G�u�BVٔl�J�>Î�Tlm��3x �p:��YUk<��~ٳ�F�/�A�_~�����2�Q�M���9$����e�-n� ����i��f<y~�kx�9`^ڎ��!�e�V�<���O�z��b�d���6��M�ʝ�AW�y���-U�����ʕ���� EUl��
������lU�W�<6�i��(��W�ܴc����]�����v�M��Fs=���wg��1�ՃZx\��I�Kal�s��)�;�D�*�6�g�-��|�����0��3E"�"d�r�9��4A6k!�M�����U ��/�Ǖ��FA�>[s�h�i�-�L��tޙޛ�s��?����.��Z8��"w���������}���e��n�Gx�І�&&����Q@B.E��$R�q?m��3ڬ̗ȳ�i��e#��q֦����I0VF�I? ���q5��咊s�J��ݛ��^���o^nn��?�P��! II���r�68�a&����Y��N���5�co#�'�ZkCwUWX�_?=)�O�ꓯ�g-	�2��˒�O�'RI�9�q�,�<�<b�y+fZ>�m�� Bv�Rq�ۀ��)�|i�<G�As/�±gV�OP��u3���#��cgx~*���ٻc���&��|�ńa������>�̙�=G�<�0�����w|���v��w�eW�.����
{�Uv��j��X5i��+�֝�,����"-S�y�|���3�WR���6[Ϧ	?���kx�7�Y��9��,n ��N9�C#��w�e{=+��Q�B���1��_F���TR���7���n9��o{t��.ם^�*�(Ф,`p&[�*A��*zy[��c7���@�q7F� jU�Ĝ)�!M�.�↞^QuYo�B\�Q�1{vZ��L9�؝]����H`=��&˅q�gN3J�E�G0J����o݆k��#(���G�6�FY�O�/�;L�N}	W����S��*^��i5��Tۀ<�`���+r�o�\���Ylv����*w���ۑ�"L�8����d���\G�j�:�}���6�,Ұ��
���Q�w��.�k�Y���DY�j������������@{d��U�'�R���3�%��$��P�D�O�w�(����A=�����{Bm�yq����F��w�N��]����k׮\2cٽ�?�N�o����c�~��Ό�r��:�� i����j���8%t	ψ^ �Y�Mz�	gJ�W��Α��Ɨ=?t�P^SV05	�6��7�F\xV���4�`� .⼢���L� ���F������O�l��E�8�MNf�yZ��p�� _�E���D�1�E9��qT�����Ŝ@8����=,տ��]��2�]�}L��`y�*����ϓ�ì��+�A��/�.���6�S6{�<+a}��1�ok�4p �k�;ZR6m�-U�9��2�W��s� Q����{�!66�qy�$��%%J6�;�|�� P�ܴ�;�^1\�bU�1�QEW\�W���4$����i�����.I耀�FC"c�<I��
X�r��|(�,��Nl��cbemq�M�u��I��^)JE#�Wg䊒���~z�TC�.i&�C���/��Ukt��������C��4E|k$&T�uN<��(N����B���;3<#�Hf3�4F���
C�P�+ޤ��[ܪ�����$\�4�ȇ/OERєK����?_+Ro$t��s2�UG�A0V[8��{C��7��~a�8Ƃ�� J�ŧ���!����N-�9�j)�RJ��-5�K�|�$��BE��˥���ޫʇ��X���7o[�2M�*���ZM�(�#T|���kd��d��f#|֮%���=d�A3�}k@��=>	��кB��t/�g��c�խw��u�� �X��^X��
P�k=S�u|�R:�Bk.�J�ɣ��3� <4�����d������Q"��7w뮫�Z��S(�E69=.c�Z9�!/ �=Ɋ!�=kɇT�Ud��n�ÝU�LK{ֳ�o
�&qR���=^��r���CԆu��D� t���&aj�����X������y�=Fߛ'b�6S���%~~�-���(zIOolb��1���׳�#?"��VMxï����O@)K�d,���,r�w��v=J�e�-�P�߅h�9(w�܆��<f�6'~��7��ku)�ڣ��S��ȇ�m��f}>�a�u�KI�9bk�b�
�=�
�M��v`´S,�����0�-��4�P�*{U7^M���}�q1��4���T��&c)��DW[F�yʭm�=�$�z�j�[(p�OɻC��O�W�~k�M��.вHh]��9��#ݨ	Ìy$�WLI6���*{�Q�8>��J�W�����������Ѐ�����`���r��._P +g$�_-T,.�����ys���G��),�3.Y�-j-|��!V�Uz)�z��4��iZ��>0!j&�)�sP^bpC�dI�`��D�Փ�:G
}.E�F
�ƛ_�a���:��</�'���jZ�U���]�eh�\�X1wv��N����p�J��ތ��|!AB2�cbrJl�F*C��ř�o�UT�@Pĉʰ��?�y��<	j�u{G@u=2l�E�`̿��,R�(�5aH��;��#y�mP��O��[%�@q]I)�|�+��S1��E?�A��ʷkcG���=�P��a[ѭf��/�l(��C��N��-�>�s�Rl|��-d�'2���4��p1�_]e�l�Œ'9���X��eL�%��Y�+p�]�����h�����ўR^���n�r� 5e��M\*�_qѝ�CT��Ã�y*9+�����qcVƿ��f@�R00�0X�6�ld�0��`+���5�]f���]�q�@� �Ǝ�1Љ��]<ůy���h����}bݠE��DO�+��	˚4���Syx��)Q���1��X1��X���2@$#"��k�_G�����F��^?̤�.���==ob)T5s�\4���]�/׵�.{�������:o�@\�A���rs���y\lq�Jh+l��8j� "��$y����͜54�ZQ���ރ���lQy��<2�;榴I�Tj�خ�91�Y'q���JF0zR ��I�<�