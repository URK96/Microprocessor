XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����x,*�hs�Ey�vmq=�t�nAO�����AG��f�L�?_�y�+RжQ��n�id�NT�
h�̐��<�8��8B�N��i���s, �2L;C�IL@v^���GY���w����Z�\�SBn *���}<=q�{l�$[p����J+�7?�̕�JqA�a���-�@� �Ć�Ä�0�Ibr��.2�����T�$Fs�����lv�,x+'�_�yN�0�<�kp��J��>��ڱo4���+"+��i]g/ᬷ]�;���=e��Oڬʭ�r�;;��,�Z�ʐ��l���;Z�����4(<�'ӹ��Os�x�{B�} �
R�q\��V�jow�"�o��*�`E���P��^�4�?x���W����䛉����F�����|C_���@�xrh��n^m�S�r>���_��4;M��tP��W�\��"�-)�N����v��.U�Q��Q�(9�br�f+���ČcV��&�x��sE5��!Ґ�9E<{ap}����d�"�/�Z��>!W�~����8mT���԰D��q�X��RӑQ���OL2e�� �JLu���8_����*�(/#�Ç����Oa�Ï:ƌ�k^q�Tt�E�W��w���L��w��K)l�a�|_RU�vذ��Al�"Ob�U����C/���$�9H|n14��(��Z�JA���Uȟb��%�Y?������I鲜;-���F{�����$I��e���f~cs�G���lc�1��%�֟XlxVHYEB    b892    1b20�i�n ��v�`8��"���1��QZ_S���"��G�����?���cƆ��K���]����R:C���6yG�}����Xz���Kם�zP�.L��ez�Ԯ-��i��SBE6q�/�Vf�BɌ/�:��AE�Q�f�����ױu g���(��-Ş���	,��3�{�إT���p
��B�҃����f��3���t�[���Կ�!���w�u�oJ\(��:Z/�Ҏ���N���:�%~ ��'�chJ �Z�v8Q �
;�p��>bj�o��	 ���ė��0��=��E���ldyڙ��}@����c��[�k+��_��v��{����b	̲Ᾱ�H�܁ܾA&&��)n��`��{��>͊޶&� �aԨ���.j��R|�iH����/�h�U�0"�5 +d���fD7b�ׯkRʊ.z����`�B2��&C�鼬s�Fa����]�9?�?J��M��Pxș�՘'B�xP��J����4|�|��
�J$�?8/�{�ɾ#ʃ��Ϊ��Ʉq�{PJd��"�m�2��K�U��Ę"���V����K�f�^}��q��:I�����ҿlhr��?����3�)h8����5[��R+P���!2̈,�l`���ˣ�G�viߣ��
��?�'TA�\?�/�F��)��{�,������=�C+4��`f�����C�n�m� ��qB\��5�]2U(���x���4�rI����e��c��PD<v�u �3�s%�oW9�#���!��ɹ�o~��gُ���6��Ax&˸�e/��e�R�~f{ԃp�Ͳ!�������WU�U�)�����Dz	)R�_�.������ϕv/=�H1��G����Xܵ��=-����̃}9�V�.`��	k~�!���Q�;SvzP��A�L&���^Exo��oE�G��]��W�Й�R���,	�;������&'�q�WT�N����޴�85��AK���%�ufZn{���»`=�1,�Ej�(��0݌S�ޖ)���6DAp$N^�1O&�aO�'	Zɞq� ��.�$�y)XSb�>����黤jac)��2���X����������z�F�~|�!-R��O�}�l̟�����Ʉ��{�ou�����[��đ�����~���|�}��DtĨ�<;|�����$H� �̤�����S��?�����4�4w��I��On؛fx��J���far9"*N%��v\�Hx�#�MU8E�u�)���F��o��b��P����+'��2u3�@��~z��	˭�.�Xz%�����U�6W��iu�l�X�����Ф�C���W%�ߊ"M��;^�	T��ƪǳ�҅lݳ�-u�e�Al�\p7�/HSK7�!K�Ñ����9�`�HG���R��[��a(�,hD�q�u�/b����}�ڷӟȇ�#D��ȣmk�?QK�lc9���ƙ6��xׯ��#s��l7�'�vѯhf3���K;f��h� N=����pry	���R���i�0<���_כ�4e�Py��������T�2-(m�nP�|+�4)�j���
�-'I���<��b��������k)�7Z���Β���X�<��[_��v9���g��*��,�D��xP�
��.�}Z�Ӄ�xu@�_M�t�����3�g�fix3��iasc&w�{���֏މ�������$���ԅů�<�n��-X�t	5�r��N��0��W4[�
a�׹�x�@�	���+�)����6�=����.��rXp����hs�.5�U��
{�t>��B gO|�*���Ӥ�HC��1s��Tܧ�I�$�\k+o
��;�g�/1�Jjai�3K���}�m�hU��r
�/W+��j���2��a?m�hC�.�r�S����Û�r-�iڟSt�y�怞H�F���uO�SH���ބr��7[�Z���
*ثӧWFo=w�c�x�@�I�t{��i�@>�3���A;���e�.�6��%��q���fd�=^��܅��f&��>jC��,�|���t����x�O�Q�����߸<S-EL�eN������`�I�սА@>��ڂ"�L;�L�~F�R�����Ѣ�_���B �jCƵt�,o�y��I1u-r���=�Rx��	&� _�|u�����w/� �lL�7��
�R����Ē���]{��Dþa�����>"#�Qr�r�h�y-5os)�0J��'����(�8KV"U1����2~4�b=�yH/�歃8U�W�������#z!F	��Y�ͯ�z�	�h.W$�;�&��м�Q��rԁ���zN�e��7�_��)�oÁ:0řSn��FG�>^�XJ�5Cfj��G�����I�,�1���Q
�C)9���sG��O*M?*�J��<D?�j�0��e
-_ʛ3�ʉ�Z���c�AU��[^�C�<��������vau�$h*��b2�!E�b��K���R�#�Z]Ң�{\���y�f}z�֋��r�'E[��!V�"��:D��'[�~��H�f�|D�]36*yC={���gO5���x3�T��@�5N �%��)�.A�K�6()7�s�I�����Yf:~\n@Kt�o�`>�y�}LGA�m%�Eg<u㸊c��e�t���WV���!b=�������^�g�A@f��!�{���U�m��;��m�I�X� D��BS�vQ�jT8t��;���uس�δ��+�`e�e̩�����k<2 ЩG�7��.?��-�	��7��;�bl}c(�n�;�f�7������ *C�����8�&6��ޖl×~5��I�Zi�5�^�u��s��:8.RKm7�� ��{�]Bӯ}-Nj���� �[N�k�杚�V��V�C�ɵBEl��H���lmǬ7Ëni.��U|GL�&'X�rYQ���[V�L�.$�r���q�}5�|���z��hA;�=�]UT����Kը��7;�r��w�_�/�9��~�����~�Q����rL^G$�SݳgJ��H�rD��oe���.d�A0�d�`�E�f�H!�i&%���9�gb���G�epl��l��Ʒx7��P�\�&�l�?�I��B�����7�3�(|+��������]�\J���ta#��@Rg�6p�����"1�*���_����>�n4�:*Pv��&�݁����/���b@��T�^�ةf���Rh
 �\!����ұsN���ս���E��`��6�tu�-�T��1��"m^Re�������+���n=�#��>��m���"�Gد�sm<���0�>�8&<��O���W�/�;m�:W\j|
�G����E�Y=M�@ʿo��ݙ7��������0YaR힩*C���v�\���F0ɱ�)�GbQW0�O�S����8�F>~:Μ���Oq*@�J���굂�>+Bpa��y7<~5W��?����Y.��4��b�ڸK�R0��j�h{bZ��*����ƀ��2�y�0��15P1W�q�y�==}$�ޑ��@����~�^bL�G{�a'qy��R켔���"B�_N?	�9��~�ӧ�M��J��(@ɹ�WE��>�cw<�UH�Y�C�4�Tᱬ*��y3�}҈6;(���)<�3v�W�\�dR��Aӷr�3~�$?��D�Rs�N-�M_�\O3۝����#�@lL�C��2T�`�>�[�l�ebt�1y/�T�̥�\��AIX(�v��g�������K>�Fv��wb��}|��9]�]۽[{]qJDW@�>+i֫_��y��%2����d�tX�O����ַUMM����Q/�����n9p,�$���_�od�A��HO�M�k��5��UT���a*�%қ6�im~��va�#�uF��Aڐ�c'���uzN�(X��fd�>�$2�i")��ʺS�0���A�C_�S�������e,�>1�0[��j�V��F%.�7�d�����W�i�J^K�{]�5�0���.'�U�7�pZ!R���
�PR�d�E������q�cͯ�Z�ߩ=���N��͠ʞ �4.'?}�So��+�������}D�$	 !�B��&en��T9�9����>�妠KO*��4t��x�%�k3Y<pc�V�r%f5 l)$��4��8)A6�u�� !(!���֖7/PW�@hvX����*�ť��'i���soIݖ,	ϵJ��J[�2�xN������9Ӷ�!ړ����I�&//V.+�J��3sΙ4�cTY��Ƚ�9E���x����^�I��$Ww
�Q�cbNQ^\�=k��dO�B�Ǣ⃇򔷱�+�-� ��$@�7¯d-�zU�2��=�s.B�x�(c�2#����mĪ�zw"���T_/D���L(���b��n���wp�`.����L]BHYcQ<Ӈ��Y#�6µZIcV�L��*�P��K�Ǽh[x����r:�GG���!�ࡹ�2[����G��g�n��@+��FԐ[��Q��^�U�8�vjnJ�(1�/����_{l�UM�r���y��V	�9S�*]��bS6Vq����ɚi���@4I��fR�ϱ�(,�NHf�^��M�23^f�,��F��/c���J��5��w���{۾�]c�:�Y<(�n0ۮA1dj�gIO��K�)�9��(���� 9O���.鉤O���$5�>�1�@�47��G���6����������� G�&$]�u���#�U��]#N�%�7�ZW�����הz5-��m�R�Ć~ �Iw� LR:�(��h
Ȃ��G}�{��u�^_^�#`�o'�rʹ~��>�\��EYR���'_����� ���,��)�ꋾ���#b�6`_t�T2�%`�[�>���f��q��n�/zx��ER�˵w�.?%9d2MK!z���������+`r+�G��8��%�fE�k"
���9��1���LY�UD���t$�M����(��4��gb��Z�����bA{��.�N�K_f�w��}��N=�i�P粳����Y�9�,t��$c�]���� ��Sf�_ߖ,�,����<K�RI�[r�[���;U,`*B�3(Q;oK�o�^�_u���m�>aZkH8�O����q�.��'&�<��K�)��۞��wS{� �V)n��� *!����!3e3svk�Hbh��|��q�H�Bl�Hn�Y���rY=k��S#��j�o'��H�{D�i�� |�5�[�WE��ܩ�B8~��atS_���J�؞>��D(���9�%{RA'��?��t�>k�.����T[����x��l#�{4��������z�u�5�i¦�FbM��o0������oS��q������nc��so���j�����h�涎��ǡ���ж�J���;�F?"o�]^���׷�ӿ� ��.����J�ݑ�m�&jk�%��͛� �U	}�u�C��5�ߛ�%K���`���=B��XԔ?e#��*o��{/KOʤ���Hd�ˣ�ߑ%h���sA�m��+����&���f(t��(�a��7~_fP�"�V�3��I�|���M<�K�w�ˆ�~0�����|�8�^X��5� �W �R?�J�E=�>:�5 2RВ�[�iNX�H�� ��Y<x��g��G�j�p���^ �1Տ�b�C�j'OrE*�~Z�Լ$!�h$���4h��Lm����(j]�.�^��&�-�m����b�0�����s,�'^�MyQ'�N��S2cyI�LT��D`��a�N�k<Y Ԧ�Z>�m��^�u�\Z�	4'�61n(=��8'xR4������8��d��oGKS<��ѸD��T<8O2�=��y�V���<�|�	^��=��G�u;�o'�����x��d�?��F~�{��@U�؆%�պr��y�+����Q=�INA���� "C�3m��qQ<y '���v�^b��2�����{]��m��kU^Ql@fR���/�*��{� <p��/�ӳ�w�oo��Yb�����tu�Kl��L���_���(X�|��&��>e�W�wSl����9U�P�=	E���2��k/Z�m%�g�Ee~8���3(3��J��T�Dt�����b���'���B�u��5,�����
���o�l�ɀ�Ƌ�\��5�	���H��$��:��j$��hĺ"�P�R��w��@�\?�q�d�~�e�9�W`�ފ����6L:�u��Z:j� �"F9��N��w���	R����ߨޯ����=9�;��r�aeR��=�M1m��N�}M��#�^/a
F\.������t��a��7~��x��(�@��L<r3�b��p<��Ȓ����gG�ih|�!�a�C�Z��547���CS���V�2�ݻ)�y�@���a��f�i풫E� -]rLQm'Ђ�QB���"�3Fv�؏�@�H�ݡ�w��Qt��5%ڙ�:c#$c�jS�Wnl�9�tZ�@Z�;�2ulJ, n���#��-���*Nlv���V����JR��>F�"k��է�uM����Nl��۔ã�wJw~��t~ �P�nsK�[��;�A�
hM����BW�*�\�%K�/LW�@��������QrC��PQ\쟭�o�@�q.�*�y�=9c����6lV0b1HC�^��wW�j������[�v�S}�A���$�Q�74�%mQ4F�\��H+��lj�:SǪd�o�F�pHΊ�$!>UFZ$��Z�ڞ%�f�J�Qm���)�#��G鏨�Ć�]�,�<��LYs���c��w���gw�`��'x�*;��خd����")IA=P/U���
