XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ҌU(���:%�
sm�("�������G�.k�C�����]���<�_��m�q#W�L�䄛������&����v�	#">)2�-�8'�SgEy�c!�5N �Eqn��	fG�鐶��#�;�f)g��h�,��[-���Ǣ�޵[�򨞘�u��[l.�I�M�~An荙.Y��ri�h*��U��=XH�@|T��$[m�9�Lwd^�/��EV�����/ߤ����'..c)$K�Vo��l��#�!��6t Ȓ�!/�$�t����K�b��\�"��(�CBAwq����2��al��U��5�c��`�r�eɏ�����|�|��^0�����r �����(�;BӉT�TV�2tZI�B��ᙩ�q��ι��S�L�Q����T��R���!M���#!i��Ih������)`� ��]J<J��آ h��J���Ҙ�i�<i�Q��]Ԭ˒k6���( + g͡G�9X��n�Y�c/h�n��܋Sݑ��c�S�����nM�*׽���4%����-h��R�}_��W|R������4X����ɾQ$	����7�1-�`���L(�zJ�#_�H�M<��E���T"��Y�ׂ�mqM����+?�o4�(/v���]�-h�-I���.:�v5zvqlF�5�ތ(��U
�=IH�y߄f�ڵ�*�EB3���9�}��D����F ¶�P-v��G�zP�-v���9�R��[7_�)_�H��5�:XlxVHYEB     b88     3c0���=�i���
��s|�'�W���0��?��O�y�u�gc͒w���#4E��7;��A��e�SU�z���.��Soՠ鬪6��x�ܣ*\�D�^n�S��H����l�x _����u��P����';.�ퟏ����J��������MZ;h;�O�B�C2��\��B��K��X�VcE���X��ƴ+N����HV��O=�Kv[�a?@3�_ G����Ɯ���ξ��xU��H�YsѺ�K��o����4C_PNo��G�^���-�"����1Cc����:�rY{�+����J���d�K��ߣ+<Y�Ի_��u�cFz�Ste����:�'7�J��֬kg2���	0��|bj��Dn՘1����&����ۘE2���X��;�xwq>	=�������,�����eRƃ� [I�4w�c�U�a"nk���W�Y�dy�?
v]�?<�2����X��w��T� J
n�7�l�Z�>f�ޘ ;�c�����N5��߁Ft��,6����#~���ݦuI�v^�d%k�ؚb�i���0Q��[?aE�m٨0���O,(��_3��4?ҙ�W�	;�N��K��Ȧ��/M=�3��ˤP�`&�o���� #�d��y�l��Vɖ��N���b 3����D�0�j��I�aHJ8��S2�bll�W��CR �d�Yc���� �v�~�V��y��˦�ɦnqg�DUH~N��pHU���wd�Ȼ�������Rf��5�T�F�#�*s���O�������Ad9b�c�N�\�����o�����7*kCH@�rDm��W-M��a�	�|Q%�S�~�k�Ǯː0L��TD�;B��d��8߂�����D��&Iy�7A4u��X��ˏ�\n rA�K�k�Z�L�O[ed3��`O�
�_����h��46�-�.ۑ#ce2��*����m�bږ��