XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~�a��y��� -��NK+~�F����2Y�EF9���G:L���9荃�J���o����9�B�M*�VT�d]� ʮ�?o��KW_�L���gZA��9t��a�%�r��9���
8�s��(��L쭶|�2�RB ����X>?�ٚ,lE���u�8|��l<��{�g���%�-�1R�	�Dֲ	6����1��IpҀ'�^�}o��� ��zW.��I��4!���g��b�����B^�����F2���t��5�p���S��/cst�5����\b��|8��j�� ;������_�"/���{�㻏���1�#��m!�wU� BHX��8�4&H1He�)�!X�.�P�F�b��qt��؆y�օ�G���!�����Z��xn�Ƥ��Z����nn<>F=C�jJ9�.J3�>1�a�Ѓgǈ����kϪ���J��Xb7�r��Nao$0_Rzo���I�P��xݰ=�f0���w
���C���	�&q����o�k`>pؕ�M%(x�M���8bN^�a �L��+��6��P��Y��C�J�2�Y����9��;� ����yÜP�O�����5���-�D~���*h[��
bl�9�]��ފ�����5�Dˡj"@W(\њ�MI���m,�Q����z�9�qʬ$����Mޤ�)�R)��J
O����Op����I$�/��8ND�3��n�_$lG�;��2�Q<w�{u���ڋXs�uG���y�:�D�Gg��ss�c�؄WG	�,XlxVHYEB    fa00    1390�*�%��en�Ԏ���8�o
�8 Cd�':$a0���g25#@c���h��bvIr>��B���<���t��R ��s�P<X�z?���v���w"��������{Bh=}�~0��4e���o"���<�}����\i+�*�t�@��$i���0àF�!:mgX4���"l���D:�9N|�w�V����I�D��lKg�޳�v5{��D��Ҥy�>�;�@?Z)��IU4	�d�
�SQs<G�����<��,7�Ǝ���>i�meE�3(��6��C� ]\��ܨ~��	yQ,�%K�Q�O��mFq�sI�".#n��lu�襺O�a7�d�k�����d���7������n���[?�u8���.��baI������(/U.g'�~�0��C��KX���ݮn�����Y?���:�4�ILlj$?�2L��E��Œ���y�7	`"����x�p�Pc��0.��w˷"QW���s�5"��V�0�JQ��o@��E$�bx�9
Ug=Eeg�ux5 ݮgD-�\��5��L���7m�Y���f�qD�CA-�b$�VL�*�)���U~�^I$
Ia�|=U��M���3"��� ���޹J��ꬅ-�v��W�5���"���얖)B��r�[��Ѻ�`a�_Xh�<UفZ�zq	����	/Ǣ�C�f��N_�noC�dxW\8Y�.d�_��
�m��H�\�Z��v����ݟmi^jѺ$��mi����GZE���Y_�p�dG��7�#�5mJj�����#�R�|nNT[�z���_%��{���̫s��Hyk�Q�! u�C���Ũ����G�Q3�a�(*­�%pD��?yc���[֣K��#`(Q�N�Nͩ?�M�M}I�Jg��q�8�����J� �\m��G �C�7	��:~�����"�7&=Z`A��A���B�bZ4
�,�q��?�B��T�1V& Q�C@�M�20:���wP!�o8c�2A.���TQG�ߍ�!C��� s�C���m���o��E��j��o�]R�U�����q�'��Fq���������Ƀ7��\��kc����H2����R.A�
+:��͠t$�h�^C����/s�?�923��*��½(�|��)�6�}9�F��m��t`�դ���f���PP,������wJ�ƹ2|We�٘m��&����KF~�曩�g���C*�g�\��))Ks���Ԇ��fL�!ꍞ{��Ȣ�$�V�[�ƺ�ݭʥ�Z�nԓ��(h�_��p� �U���{����.�>�
�pzS?"CqM)���N��=)j�K'���:�ހ�`����[����Ƌr�9k-Y�::i���϶*W���B�M�ڐ'��B���az*$�������ϻ(�o���\U�W��C
Pw����v5cz֔o@�_��j�T)G����+��%N{|�z�&}��3�H������_d��n�e��?�����Z���5J�7�8r'�w��l���c�{`�_gE#�+�4��W����������ao+c���
d�f<�d+O3.����X ����Kͻ��CY��o}!m\�*�" �lDY"�5J�����~�S�Ȥ�`3�����r�CۀDk<�ާ�I#uu��)��b|A���_�M8|xi&Q�UZt�-f�g I����
tf4t�����K�F&�&t�W�AŮ���[�CB�V$jr�W�����D��i^]魰����"��2�c�ee��ְ�r�Su62آ�Ĭ�7�l�4��5{G���+���5x�,~�f�cu�%�Lן8Φv�F5��d���Zl��(�k��������h'�9�<��u���S�֜�K�"�LD!I�-^/��8X@=�ۅE~cGx:1�V-<k?�x�G��4O���Q�e�C�!d�&�sd޺85eE�ct�{�3_蝱�9m�;�Aw���<�l�ɧ�_j��kj����T؈�Smok��m��|�m}{��$��=��h�d��t�Z�|�]��˦c��ϓr\=o9f� �H3��J~g�I��w1�C3����X{}��|�A+��� �������7��2~9ۯhF����x��,z�>��BG$�l��^e
�;E3b<�K��I�{��7�g��=����,f4	��(�@��M�������3>�5-�^3�g��	`+ACE��	��V�Fk�� ����!���[	ȱ�c��Oe��i��6�ԕ�&`̋l4l»v3#����fK_탿0)�L3u
�6��J��``!߭F��/y��o��
G���OpTIG�iǴ�B�A�w4�D���/H#��#�N��p�<C=�f���k�Y�d���@����$�_�ێ��߂Q����mX16^��+o�p'�0E�;�Z����KAt�p�z% �0�����l���R Y��6��[X֨ZH?ʏ���
n�Lb8��ߌz�kH?��H�	�jlM��,��y=_���oE�0v�e��/�ܯ���$�mzuV-��4�s�*�xZx��=F�&�w�,\X��x�k(��{j�N�L���V�:��	cB�jw7,uڼv\��
��A�8~i��&�?�f[��$#2�{3|��^-�m	
�UlY���\P�4|eл�NKv_](����A=���|�[e�(�w��gq�e/�Bk]z̘e0�4�_e�P�DYJ�c_��"s���q��ĉ~k䇗:�E��}C��QU�}���U�b����0�΋xPzA��:�_���?�T�����A��J6v���������>�i��d�r!t��Ad�O䧻!�d���Ox���ᚼ��G�����LdZ�<�������=�|��[�����s�����-�%g#���k�� ��*$��= �>���t5�݅���UWD�y�!��r�7�_�G���r�,I5(O�>�s�Z?����6H�vL[�f:Z
]����	�JO*�hPI��wg�&\R*U���n���|�i�/��?4��,�[VJ�iU��a�42=����˰�z��/ր8�Z�vWi.��k��&��Y�
�&N�Mx��|2�!�7^]?�i��1�lh�ʉ�J��ᶤ��K��]���1-6�LH�]#]��*�X�����R������}���3h�J�,�n�6x/�ǫ�e.+-`����u���E�������
��*�A����Q�T����,E����0�f*'~҉M���ϐ��!���h�I�6�d���|���E�Z��ל3�=᪎'Ү��Q�-�饔��N8o�b6u@ޑ�|���k���bf*�v�wq�$��2O�dN�ێ�9���^P��d�wڻ|ځ���u���\�M��^2��C�uD��X��x��0��y�O%��85����Pv�v%9Ȅ���t�~&����Z�g8?��݄����P�
z}���ț7�D�LV؜��Z-��w�P�+jӲ��=�?T�Mk�g�Ww�?J�"&b����|�.��K�m�e�@���	�lp/����W�>�����r�������[�9p']��S2Ћ�1Y�����"}a;!%���K�w�%��0�a����!5�w��,h{��u�q�=W��+˷�ڿ�8��w�M.]}Eeg��&ϯ��^\���� np�~8/��=�J>������5X���'��	T������F�u�M��*b�ؖd�#	+�
`���k�S��Ym�{�6@���00h�G�-՗Y+�U����b�؂�3���{��qj\��RD\��?��If_
�,�w��oE���ʽS>Zv�#�Џ��}Y�x*q�a?�R�{(m���c3���ډ�M\�f�;��cE�U�F+��Tp��{2�$Ūk!X~����ɲ!��ԘTV4w!J���8?��T�0��N�Db4�4�Ȃ�ũ��:��+ �lB��d�#mS�VY���,��B�˔�qT"�D�+�A�Z��X$�?aqvǯ'���Y�ހ����h�/EW��үoSt=5��!�6���Q���wg-���0�>�"8�ڀ�;8S���coo]*��J�N\mFA�l��F�j��g�W�I�D2< ��iO��m^�����Zq����p��_����W��;�ob2#5����v�v�h�b���>�_f�3E���CR�W'C��:��rXtʬ@�������R��2����z#�����|�*�]�i�����;��3��*X<�g�+�,�X��T�5it��Xh\�I+ys����327��޵tר2�u���r?C�|�u���o���p��!�2��E��#S�S���CfzjI+��e�e�y������/���b�Y�t ����G�T�?���`0��������:Z��msBI~Vƃ��.q�A��팑���b`JE�T��Ux�60�A���`=�A�� ��&�{���*֝��m�	DH�_�#:���nިҥ���h:t.�?���Mձ(�������li))�tM-��5@R?����)�YU��bh�u������9�M� \�_f�P�%Q�d��ѝC����7s�4���e��(6���ç�Ǐ��w�˵31������B��@9�-�Z���t�o
b"����x���[舳)s)Π�<�MS�sڠ(K��<�; ���#����@�䴄�^�M�h�9�6�.9��z�e�EJxΉ�2��o.���_'3�k��N/��Y���M!O\'��υ���7cS]y�m���ǉ +�^�o�o%P0����x ��S�201�]�;��:�,�7�j�o�cZ`T���~����o���{�K�K����&|�Fs���Y2-Z�8�1��(P��[�:Gʸb�{M��h���Z3�X�1�D�#~��{���>m��XlxVHYEB    1193     3e0,�#��İ
`�K��� ����oS�/6���@��pgc�׍[qI�7���V�7\�!�X*��,,�rp�*y#=Pш���$[Zwy�B�Я�R/��Nq�U2�بe�D���C�HW��ʔ��9�^�^��*5N�,p�D5*�pF�>6���إ2D��)�Z��6��I�ـuI�隇�M�"���D�M�'�y���,m��cB�)�H�|9Ay%��<)I&�_S���S���<�K���`y��Tj���K�-�)Y8uα�|_�Ha��.v@8�'?��iV��#�E�� ^o�W.���+�li W�Hr#̟Xi���s��(�$j���C6��ވ<J�,t̘5�5m�����Bm����\���O���Cf�`����;�9a&#|�<b�
������~�`�� �2�vL���D�߯~d���ڼ�9F}��yrL���aإ��`:@��7��$l�q��ċ�$��M����V��@�	x�K�搜�F�e3-*�MGs�;\���%Ϻ�m4��1�s�?�o*`ĥR���k�w�e���Q�O^-�-PɦzWr�e�0�<aP�Ga�Gkѱq?2YM)���c5X��U�6�W4��4��G^���P��H��;�hp�zGz/�e��"!/�ڝ]-hm���렠�[=�bE4�ZH>�t^B���4m�9���U�K�`��Ƕ#���Ð�2GL,v�&��V���W�eI��{���3�2�dj�]�p��V�nE�5`&���B�~�GBC�����=��K�Hiع_A:�-}��5���0R>:�+�����Z��K/����e��wj�d}k|81n6�#l�<f�M�W+Y�Ƨ� �ݒݠ�`�
�K�,��D{e���+���T�*]�&dzL��e3e�G�6��|l&�io�j�>���XUդ-�����GC�*��nL�9Gnܥ�ӱ�·8^�=)L���!Ӛ5��T��2��?>�C��u�