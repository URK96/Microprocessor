XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��d��Ռ?�E�C9�B}��{.��&F.1��n d�r���p8��I��>�K�}��4�����%*h�=��P��j�om��0\e�PAz�������IY1�����1È����}�-	$�.3s:�q��VJ|����j^*L?�Ї��m^�ᷕ�-��:q�@� �:0H���ؐF�����"�:)]>0�?��b/ Q�Y�֑ǗQ�饷���1�}߯֠�d���(��E4S(a@	i1A�t��L�昱WX�s�/uj�y
���^GL�ƌT�*P���P�FɛH���2b�d�=��9kdJ񨣔�z��
z%��B՚�7�}����C��{���/����+���r��\������)�b�]�^���p!�<��)���Y���������zf���l��ؗ�D���Pa[�����w���� _J�Z~�b�!Ӫ����� a���5�� ��uWF�XN�0%g FШR�A�� �s6f
z#�͊�4q�`k���^_�O�ū/LE�s�YP�x�>�E���T+�[$��;s�?�WK±�1�����m%��-�J^�q�I�@�˫K!�	��N��*X]�#���c��ԓ9�ܮ�~��4k�dI��	�D3	�-�2��?�A����5���"tU����|�׀%�[KL��h����߲\�lC�U�>��z@�D$KV#��un��	Ч_m���>q�Mt#�Y8*f���e��{�-K�F��3��۾'����b,��̢�u>�aXlxVHYEB    2b30     a30����Kp$�c��9��\�:���� ^�
��@��T���a�$�F$��gSbC5w"G7���o<�y�q����n�L啘�	Q���V�m[֤)̸��]s�O!۫_�.q�)Ty��4�Cn ����5���Pv�
2�C����� �$�5���,Z�<id�h�!�N>TTn	3�E����3���:FeǙ�2�D�p���n��j�i�nȮ����c��dV�s!GPE�Ҹ�:��ʲ��l�INv�����J�zT^L��N�n}��	�E�� ��:��>�x#gYv�C��\N���?�S6��E��5���[:���r��u��D�&��m��n��2����:��B<����Z�W��ou�������w��S'���r��#L��B��9�^��1�6Q1n'�l0��U��Yo�{���75��_)vF�%�u5��}ܝ����ט��t>s��,�o�dSa�1N�������	���c�"畈R�� v �*���	�Kܣ���7VD�NB`>�U��C"l��t��nY*��!#�N��gJ����<���dq`�&7����-��3o;�P�����t������m�K�_��O�K�x6��J8�}	7��>�]^� R�õ�әH��M?�Dj��vf௺@���.h�n�Hw.�㧋.��p+��O��ׄ3�-m��*�Kg��ܙ�BoT�I��#h�
���^K	L$��E����
J �j^�dQ��r}�����q���E�v�*!}Q��"��r! ����:�]�ya���,��N���t��B��b�2��� �a|�@O�����`�d�B��?'�������[ˑ�xBA5��Ji<Kx�q(�t�jϹ��)��q�TA��a�%n��+E��TS������D���<�?%��	õvun�f�X���@n�p�{2��4?��w�!����"W�Ζ�GRcT(�$�B���P���]_����oH>�P7%�m4�����8�F��ga��F�R	�6���^Y�k���s��F#�S��r�	.
�V��v|��M&WQc�:S�R��~l�ZV1��69f�t�" �9�����Lؘ��T���F��1�-��َ�a��C��بN�/�rK�0�%�[�;T�@AER9q�T4�Ke>�߲�����i����E?��Df���{?[��uW=(�Q��TLNt�-�0�f
�����')4]������){���~�D�v���	�U�;L2�����9% !�B�g���ww��И���+��:����8S4�ؗ� j,-r��������}�A��H�
�Hu�z<�����){�_}g�����0s,���X���:�]�`�>�a|C�3���,�*CB]i�;�)F�a@��X���g�r�H��5h��� ֌�,=�k�ϗ�Pp!䎹f�8��k��_�2�3_��g!���?ý#1f�mkK����L�)K�|�RY�R12M)6�2��J�-b�Ty;.;d�6l *`���bH�G6Ŵ�s�f�iowt��?|���K��BP=��V "�m���W���؄���փ#~�nB�gH^cFɉ����<Ê���|X0�%,b�0�d��,�[��y�L��O9�k�f%��֧�^���49�����9��K%�Hq�㼮.B�������i�Hu;����Q��:8l�{���%@I�͓��b~8o5&�)��.@/EZ5�R_ڻ�Ml�L�_�_!Vl̶�T�u�O��Q��=<�UIB�	o�؏2�]]�M�fO��}�n�U��e�NAy!��6��{�!���d.���2'����vq��/䦈}�(��o�&Nd�
pV�Y�g똧٨[X�R6j��~�]����SC�y����9s/0��X��g�5/�M�gܶ#,���s=��[��X�zV|��*$Tȗ��e?�����t��+ �������~��}EA���uB��=� ��څݡ�y��7�tF����my����j��E��)Ϡ�fRvF�/�2 ���lE890�v�K���r1���M��XR���2����[�۩����+�zWv�N�lִ���"��q�z�,~��j�Qc�͐��^��x�H>vg�Ժ�Q�%:mХ�sr�ۚ	*F�pZ��[���B}�ǿ��{!��!�,�-cW'6i�F�r.&�E0W��M[�l��m/h� vCN��=��QѸ���б��:4�_r�n�*��ÂU  �:0*8���Jr-`H5�����V!�����Ĝ��'J�"bNj�����	8�уG��؎�4&/=����[e��S� ��R��{�g��"#2U4�=(��FB�_��3����������-�����/bPr���,=J�k"��� I���M�{�S	0�R{��ģZ�q�mӭ��Ur��9�%�|�Ԙ��@�^u�A����7��4��ۮ��V{��x/J����j�Ƥ�ׅ���4K�MW�)�>qk/T|����;�х��j|RM�[��}����Y�pMRܝ�5*K�� �9R/��M�"��Ytw��8��r��0�,�{2�CoN�e���/�����V �A4����