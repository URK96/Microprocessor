XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����)	��#�#.�N�D���R�u���b�>���,����81I����9��	� ��ީ̀���P�B�t�=�-������^2j+\b`��ф���qO%�����A��i+�6$�����.*��(�7��ll�Ow��
������;��Ӂ>�ϩ�8DL��O�Ϙ�W�J�zH9p�1?�%�^��L9(�yۚ�4I0*�q���j����ޖ k+S�7J�'�?aq$�v��Ku0;�+���]�>B���,I�Jb�X"��RI2:�5����
G�K,\��{�E����[��v�L�K4iL�RD��	`��\�,)��G�f*�n���I7���+��]-��4w���6��G_��M�~��x���E J�Z�@9��9R��0�ͳ��h��x�G瀅�C�#x���ޘ+�0߾���M^�L��K����,*��Mۡsw5#F�h����9r�b#R�;"�\Y[~n�9�<w����X&����f��������vQ��Y�S-=mJz��'V��O���r��Bs4�,4��)T�Pk���g;�ގh��U�=�p��=�Ki#	��q�wW-��-C�0f�"ۃ��ꍤ�f�?R��ʜ�&8@<�k�;��5�J��*��	�>#N�j�������6���pG����;�h�,Nڙ
�������wX����i�2�J�s����B9������0��(�� u=]��YXN�U�0=��XlxVHYEB    6fd8     c30�(u֠�=�i�ܣ���7���ݴ����ݹ�U��q�͎i�F
�I�9��!��+K>����5�.�E�e.7L�X�L��@���Ҵ]/�����{�Ŝ����<n� ��NWo[��k����Td�V�0������my���p��0Y&�r`����yc��p���q���zQ�Y��Za(��<�)&�Eӹ1
�QD�o�x��J�n����i=����p�m{d����Σ9dLZX�`���j'@�ج1txi�Hƥ�M ���� r�pdsn8oC�8���ƓX�qMS�&#h+0a_�|��m���Ã<�Z��fs?�e:m&<��N���5���FG�ȁw0�Uݨ�]
����i�T�5댼U}m��[7?��q�����Fą�>��Cth.��u@�O*5Ml�:�1��G'�j�#c����zG��c<��� F���v����8%�n���K7���O�g��pG�����un��S�}���l�"KWwL��
�'U�݊m	�M�P���;�RO{��m�;G���ap��L��E���ы��ls��^���$�j�w�{CK�Z��+�R�ȸ%H4���8�����Y"�*pƄ�B,0e��<��)������&@=�e�}�i�j�=��R����".��-2upu:������U�F���uL��2J�i!�C�5���	\�w
'Z^��Ȑ�.;ҏN,����#�'x���`P�kr����A�DW�`�L�r��c�N�Z�)`�g�Ӗ���#�bޟe�F�#���O��:�1Dw
��P�I�@��n>���z����@:Q���/�C^�cW��mt��mO�;9��M��`$���2C}\)x�\z�>�>�"j7�M'������j�̸�wbCZ���xcm�*��QXj�i�sl�ŉ�����ؼQ$[��Ŀ!7�/�����uv��<xH�����Ύ�3Nq"��)D�/�m��ǶΤ�_S߅ Cfx�1�B8�dq���S�˒�P�n_#v�UѡkJl��}tGǒ�!E�r�b���� ���z<5��n�A�6�h�d<�3 O�U���D����q�˘gA{��5SG:KL'-�wb�\�M\77�獤���֤���F��O�!O���� ���c�s�5�l����gچ���t��-Ƹ<��r�$�Cڴ���XO�����	��YN�Uy�wF�X�ؾ���䣆�׈���Eca��+�T���Z�]w�Y��rtG:�h��Tv-��m�o}ǧ��#�G�߾l;����s��=�$M�՗.�����1�0�a-z�E�^pv`m�ⷰ$
�ݪ���щ�Fd�R��Or�b}W�Q;���ϯ��L���ֲ{m�>��[��`3RK�k͆�<�q`q̟VB��J��qu$'s&�ݸ��C�C �����5'	��9n���%,��&��g��-�BS��h
$뢥F�{�T���y��`|�"'�V�J�ǻ���'p�^]�	BH���ʣ��x��=7��{@:m�K���G�(+)�P.�^��x�ش��L\u1|���v���D��ٸ&I�nո*��/4�m�9!.�����9Lr�sH��#�*N����g��C��H<5I�Y�{�[x���S�%n��ȷ��_�>z�BjJi��V#�hC�~��@\<��-�����*�ov[tº���>�Qʈ!a��"&���\>�����\?���T�8P�7�<~�h��I��Q����b����Al#cL�Me+�� Ne�7:�e$P�M�����.��n�u/M�3���"R����s��K�DL5U	ZJ���׍�ȸ�V��4���*��'��RnU����X;�Dێ�a\l4{�&1�M7�q��g�	|�m$��Ѷ�Mҗzf>�(�ޭ�'�#�Q)��-$�x`���k�~���Y�A��GA�0�YFؠb]��~A>G��>zFl�w.P�g4e�r׊W/�����$b�VWcf/O��߻]k�	ꯞQ���/�dm%3p��W� Z+���ӆe������j���ôj�3��<&�/�xg��6X��#�BX�sݭJ���(�9��>�c$��ܯ��0i�' MfC^Um�BRoݨm�q�)�{����xmA�B>�t��K�p~FWDa��-l8vʍ4X�)#�0?~�b�N�t>������;�?1)+����;��
���S�OngF���d�c�:v��|j�����p�d��g�Ɲ<S���͡�g����ȣ��|�V�s�h1������L�u�*w���։i�������i�3��Db�m�9�G��x�T���Ö���5f¤p�����(Q�u����jdT ���X���Wr������Bnc]cgGN�=�<%-��}��A@�MG�$����쳃� c'1���^�j�3Ia`��_|��F^D�K�u�.�����-+6lVAH:)��w���Q�
т����ӨZ\�0��%䯐U�A�
3����Yt] �(�w��6q�.j��9�I�2��c��)�CKl���b��ރ��%U�� �X��[s<,'@b*�!x]�J�,QA�.R ����;�R���Jo�� oZ��Yn#C����1Ŗ6Vm��C&����'�-�`��n���D��_n����)(:�0y;�m��	C����9�����aQ��!M��3�F���q'�3��mT��ȫE~��NՓ4�Ȫ$c����ͧ.Gh�����������Ԉ�:���pq<Ra�@5�Qb# ��>��￿H�i�`r���R���Ty�jz���C�NAҋՆ�+C3����M�~˥|�su3�-�YH�Juk���� �t�إ-.☻���x/,���ԡW����Wh��p_�2|���u�f d|�q�s��JBF��vW���l�6+L���@*�.�Uh]��'X�*���)y>X�edp(��=j�h_��9uO�:�r`��I��HQ�aZ�=֨��&<��
G�F:�)9*�A�0�Dg1�t�4Ю;@�f� 1H.O\������