XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\������̋��ű�u̡+ҡs��j�5L�C�����(q'~��Z4������o��^3�.��\���5�R��m
�B���a��|=�rA%�7�v�5�r��$r�,кB{��	܏��Z��3t��r�sAM���`嵬�a�3Oջ?����n������/��+.��������f��4U�kn��4Z
��̳5�Ƶ�X"��:�5�4|�ZLܲA@@�ԜL�y�XC����G���8��b]�#�D8����+����ƿ�!Z8��!�"H8D�)6�z��+�|zRj��3���%�'r��i�n��p��S�4�$�/�V3�$S�7�(���-T�v�ﹴ��{�x�;1���T�K@�y�a�<С��?^$��4��
y6���P��.�T�qź���MBI<��6Bw�FΞ*Y������ꍹO�����>��(�(ŗ�e!�o���b������>m&�"���>����us��e����H���Ok�4��?g�'0���m���
|�k�b�{��R��,�Z}�x�U'U��ć2V��1A�x�	�	��3��P�j�Z��		���Ȋ��s��T�ŶW�SЫ�N���*��?����a� �3�n�K]V��l�g�B^adrN�|���M��A!�׭�b�S2&\��p��6Z�x2�yo��{a�R�ռ��������> �q��=��'�������st��Wf�mb��pK��#�oi]R�A }���G�ut^��� a�XlxVHYEB     b7b     470�x�1��S4��'���OX9�2ὺ�b��y��N��J|ϱƮ�@vϠ�<�Z�����b-�Q��5{��7�o�����?2�Q,���̚�N�^�!���q>�Q�����|e�\	Ȗ�H묲�{9�z4��.jm,6Y�0����祁F�Pm����"�l�ǖ�R�U*f\�I�~ՒGlR�Q����K�b۝�^x	���Z'$�}1<�� Z>�?R��|�|���U��cm[�.)��J��z�5߆!�SAeL�2|K��l�e���C�VJYѦ���$HA�h�+�����1Lիϳ\�,��o�˶��VP�`R�NFlk�G�͠μ�[sgCD�#�@bs@�O
-��d��K��v��t��M&"�On n�K��(������?6�x|z��z��  y�X���3ڷN)͋(d.��	�%*����TI�\�_e���Uy��)�_ݟ�ƱK:b�\�^���`]���Vuxj�/L���!t������S�d��~��{'[
n��_�\���X7,�U���I(,ߟd��T����[i�H�O��� ���J�o�ݶ�km��b�p����1�����=d���-$���=s�D���(\�@4�v���]�3@��ާ���fPH}�,�C�"ӟ�AShv1��͓ƀk�r�%��scH�l^��JX���?%��H+��Ԧ�Ϸ��2���n�i������I���fMB^�yW��_�N �u�Lt0�}�4֙��k4����1������|�FΟH����:9_8�����������0�2�MY?��K�T/E�Nh������:��� Ng���qB%T���iΆ� �}e!0 `v;۱���l���d�ǀ��SD��)�h5���~�M�>D~��W'z̺r����#���3Q�)�@D��5���ũ����U���}Y>l+>ʯ�u 탹K7�ѷ�\�:vv��{��\G"z����-Q�:;pT����GF��2����/ӫ�HJbM}�G�[�:2Jd���Sڑ�C ��������t�����<�,8mD"})b��9�w�$[�=��g�_��ϛ��ԿȚQcM�gS���Pn�|`Ŏ!#�tcG� 