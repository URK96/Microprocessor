XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>�����sOʖ������Х��2�Y �l!��4/��8���ȍ����K��m��Wu��m���[�M��o����s �Z��؂ӡ������LA�b;�'�"�;H�m���~,�HVu?,ĳ�Z���b�;�ӌ����� �u$>E+�]`xۡt�����kT��GZ���P#N�v��:˕ ������?�z�F�9�H-a���%y!�]G�H�N���rp�g�/�E)�u�D�6�Ha2.�`�d1ERN��-��%���0���H��$��o�z���"�5�P�|�T�7���eY*���{g�G��W@6oM-2�:�A��nڸlA�L$�ߩwUK��r�A��!�`,E�f�!�m ���U��*�?�%�?����UFu!tn�ϯ�Qw��t���2E�)Sj�8n�h�����t���q�$�����|���wՏ�(�!1��{����43@�B/�Ȟ�}���"�`��'�S�㸭�ݘK�L����$o
��`_�Ixi��x��{B�?>��!b�Wګ�2o�C�X3�����D���tӀ��Iú���J,>��5�m
�*L��;����m�2�Y>�\�x�kL�0o9��x�Q`������ę�~6�ޥ�㣣��;�=s19�
���)����h#z0�@�qA9n�Jc�_�M��G1��U\��B�ֻT��9A(����t�{E��U�o�ť]���9XlxVHYEB    5ff1    1040H�k�u�q;Fx��Ub�q@X�Z��P�����Q�c���w�y������ȷ�Y'��i�[j��v� ����Q�����e TG��w���5�Z&�ut�KEKys|��V�z�KךIy�ƨ��4P��S��e`;.�k-�4�g��Y���c����ZW!Ѯ?PJ��Z�w�yӏb�:j��܈>��
<��<��0~��.�|�C�>�+�C��9��Ǉ��	�IQL��P��y��{g�(���D�`Mm�`x6��YQdW@�s�oӰb�D��#3��E�7�f���A���L�/��N�@g�����#��@����lƩ�Hm�*{�>q�ll�T�}:v�E�_�L�k�y�:�����>��R�V�MȦ���~ء�L�k���a_^�"y.�m�3:�J�1O�TJu���Q�s��όP�竗@E�Z����=���n�摇L,��c��&g�"6ce4N�,�'w~��4��Й���^�Ò����3[�8`TF�����R��R��C������/5`�
٬�P�ՙ�G���cJ���Q�nI��܉���U}���eҋ?ub��w���h��7 �	�����w{�&���@@�}.R�m��d�C��*R�4	�������1����>��Ɇ�C�)�CZ��Rߙ�+T�B��X���m)�[=4t��&�ͱ=�|��F�</� 'V�l�/��
!"q�`<�UK�mv6*6�	.�����z��E�]&&�1ᖁ������U�p`�`�#�&��рb�>}���m���܉R�^.WM����8G�mLH4.]n�9�	F�n��Iz�B��-�۬�Q&�_���]��h�0�;}�p��\��3+R��mGn��X���t�p~{��)�����>#w�6Po��;� iI@f��*��a�v�y���:
����fS�v�v��)�
��8p�����^S*��U�ؔ�j-�ͯ��J9�*�h
�_a����H��_�_nH���y�G�C�kZ�o�7P�!�:{#�Y����pb+��T��v#���\[�M߱��y�2j�����9�c��c\��̨i�7���W5�V`�\�V���<?�NN}���˂��!�0�30/�m��x/AG��$��1�N����3�_�:D����H/�iw�m,�ߑ�A���a]3��ϔ��X����ܹ_N}���x�>�>�!=�ݖ�o����øU$�'%	I����Ȍ�.ǿ�G�rqJ��h3-����ù#yvR�{���V���AB��I��s�}����8JW ��=��Z$��?����6���CN�9����M�}V��T�{�+���>*�=l�^��,���i3���<���I����?�T�/ėv��)���6�C�z��o䥭sV2T>" ��b�#pS��Z=�k��N.i�x�.���p���
�U��Hm���6zmZj0U$/~]w.�>��V���sO\������i,�6d� ���j����(�N�7�t�f_~ �6��WF��b����;c�8�t�-B�Z�j�]��5�����T�R0�p [#�=Sl;��0�+g@z���PZF���3<���Ƒ�/����c9JJ��9�c�RF���u��"0�����N�*�L+;19��
�c�/5�{�9������2W� ����{�{[�廽���K�N�2f*�l�%2������ic[��쾨aB���'�r�Q��ׂ�Vϲ� ���Ԁ�b<����V���d w�~7s�H\G����$��v�P����2!6%}3Ñ,��(��	��)���|�G�k�E��� o���Y�J��j����F4�'�G�{�k�=�4,�N1�����׬0�� |����Ld�?5����v�{[��<jʆ�Si�k��5at{��S�x=@M��o]mɼ|�EѢ��O��f��n�9a�$��8 ���*������,�y��-�� �4	4J� ��]#�ϛ۟t�x�
�-[�˞Z�Z�"�.V���V��!��,�uҐ��^�i���r��J.{l���_,kY~��g�--#�s����.�cP�+>S�}�Ҟ�d��W�j�ԟ	N?2��q5ڛ$��)���u�9����H� ��3���h{g4y�7-FJ�(��_֦J,^��k�5�MӰ�=;ԅ�����Q�J�@����<A��YPUaXE�7��S?Lo�TB^n�V��@Ѯ��{���ό��FD�������d4RuMˏO�UJi� GkO�Kf����uei�X��m�8,�"����f��ͫ�7�ʲ���;���ڟkqYM|^5��N���,�m�3�Czw�n��df����@�{�`t���pʭ�*�1-�� ��6����V��[���E1Ċz��HdT�y�{�qk�M���~��^{o@%r����ى��	��_r讛^��b%<�m5XT����_J�.*�9��K�p7��_|��C�4�T�(.�;&{�儉49\�d�>� �1��2�x)VKq۝�4�/[�"��%\��+�n�Мٯ;�����A���w��A����*��B�2�*[�2���ur�p\�.���A8d0�9�����@rN�VK�C�3F�t��>L���8����P����$��A�4w�.j'�	���HO��C��6����_@���~�Z�^%M��6$�Y�����Y�yE�W�Ae����osvYz^�
�bD�O`��s7��E�#e����#|�FaV��Kf�m	� ^����0ǓZ�K�p�r��^_3���d+Ģ�v�x����B�v���u��da��!�X(sGL5�&��t�0a��ڏ��n�4JK`�}kR���.B��w��6[;gV��3A���Ә�f�G=�z��Aal>������E�A/����������n��rl�R�ݦ���N�@��R~���#
��Ły:��!_��i�:��	
G�k�s��6�sEz� �q�1/�5/���Z{�g*xK �f�lNO�l|�3�ͥﬦ}<8�k&M�V��"�;��r�C�SB�O���;���������������t��p7�n��j��`b�D�����0C��I�g�V����4�y�3�v��r�֍U�x��	}Ǽ�5��=],�����n���@o�ru��Uph�/���#�^ɧ��p
�]��
�`�6	Tb�3I8���z��<���?=H�X��`�����6�?Z�Q�j�r����aƺY/G��95���N7�����ұs^�����k>	���raT;�{��{.b�2����
|��z+ރ���T��}]zW��0��`�L	�[� ~��nӌ�-�#e��9W���u�Y�o�ǯ����zN-\A�,J�9E[{,J,�spiM_���f��C��6�G��V�H��?u��`��76p�P���N��R��I8�H�����+m���� d��*����Ww�__
V@�}�)�2c~ U+��K��!��KJ���Q�H���r�U��&_�
��=j�B�Րf�JCR𫼋��<�������Z�w`D�%�����1��
�g��� q7٢~h�W�A�5OrxK���)����-�.���1��3C��:�*�<qnP�$j�H��������YB�2'�X���꫅K���Q[�B�j���Y�\~���ʽM�]e�b�E>���~�!��:�ç�fל����:��W=-�V��آ	;�b���:0e2�$6�̬9�`J��̹K�6.Z�����0F;Y���������%���q�1�	2���x���z�xN$��,cI4����^v�������Z����P�D�>vq����7d�J<��6�ѽ�@"��\�'�O�[��Up�hfn���KQ2&ޮu��3��5�R�d�(����\�=d�-0��K��xxDZh��a1
Ӯ�p���Z#����4�ο1p��F�/�5F�B7w7Ijr%�^��M��OQ��hukLC�-�b��H���5Ʃؗ���i,ƟMkEP1��Z�2����*�&ӁN�q��>�Ź��fiy�.i��$A�(��