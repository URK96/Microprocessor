XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����r�p�؃����ʆh R˚�u�t3�@�nr����Q:ݚݤӌ2��27�����Ь�+xg� ̩XC�˟���3�9"�����I�йm.�o}�9!$�����m��Җ���Z�z6"C�{2Я�&�)vgCy�.rr"3&58s1�t�*c߫җ�t�g���;c^�<����<���a/��s������h˹��E}�V��N���9�������k���y
�/S���ڶ��C���G�ITL�V�`L~p�SLg�x�Uo<q)���Ey�Q+� �Jc���ۆU"�{�\���&�!�E[��l��V�Ir]�F�K�m�]�r,�r^�V�c/mr'�g���K�r0�/ߏ�� <��P+��
��?�M���w9'�R~R`V� pv2�~@�3�j��|Ն���yGN���ܢ�@�b6�t��
� ��Zn9�"B՝! ����yh��'�v�I��5?�aa�??҄�La����0�@O�DF��/&�L��]�=���06��B�E4�Ti<�sD�hv��*��֋j$���	�9������}hֿ�B���.������.�F ��fNф�-�i�qg�6�3˾�4:�-� �\���R�����j+	T�X>���$[�.(m�����*(x;���v����Y�TF�&�?m��q�_�lN�f|JQ*yd5�4�4[c9�|ب관l�^.ˬ���;��$'�G�b����=]�x��Um��"��;�T�B���6�XlxVHYEB    1cf8     790� D� ��惶�3�~@�&P=�\���K�k��c�/�L ĺK�"GL�t4ëXLxF��8�T�@Dόk�1���2����f��+��v6����;IE�$�Se�K�LNu(������ %2!Ϭra vW��B�Ҋ���(�r*x�o�?��}q���H������YRȪ� 0�E,=��µZ����܊mؼ�[�����I����t��G�ې%���9�}R�7G�s0l��@,h"�{����82q魎aE?�湙�WLt$^`���F!q����U�ɰۤ�D)2\Hsc���Vb���aZr+6���n�v~�9���%;�1��]	��U~��aa�p���H4Upw� ]'�ѓ5�Q�a;4X����\F�׉��%�tOy�X��A��]TM�G����2�V�����&�;y�n�f�Z�؇h�-�$n���7ڋS��x��GR¡_������)+��G��P�Q� i7��웢of�T��fe���a�n"%J"�����)�4e���_r9_(��٬A�H+L�np*�ᇦ����һU�jӅJ�C�S٪�3�� ��.[	��15؄O�+~�����5�9�"�0P�8�"���@����ۄ���5��&��U���/��'��QȘ�#�*�T+�v�-_��H���7�/&n��o|��?�;kК��V��R����kj�'I���'V�?�|F4��E��T���Dd���M�5�?p��|N��n����Xͯ�*���^�j�5ӖV��+@b�N�]����B��2��tؚ��YT�4reI��q��y��H�=�p���U%����n)���8��Z�p�Z�����Ϭf��ºc_.�oՃ����O��ӥMQޣ��@��Z~r�ņ�Bt���&�.�9����@�z����]�҉H�jC�n�eVT��\ޤe���;c�9���Liؾ~�fO�f�(�r��&XaX<����~KL��6��;�8@����	q��ߠ.;�V	�j��k�3"�#��g�N;�mW [�0hirm^0w�!j�,Q���G[�ݼ�23�+t�[�$��.�p?	�"O�&� R�+G+�E7�$@��G[�I,�'I����a�t�%j-���A�Ij�OE:|�:N�~)UʂMȰ�n��z��Z�<�?��xZ|��U� ��4x̃Z��g۷��W���~���4<�H_�S�^~2��X5Ai��,-�X5X
)�\�8���</R�t̖� �l��7�/$���<0��� ���8�q�ah���J,���kH�O�걡z�ZӰa�������E笰�	��[�ʈO���� ��Ph��
%�VP{�X':�����rI�Ļt����� �#��� 2%��2���S���������"�L���
z��1�ֿ�sBƄ�8�ygE��G�Iq�;'δ�I�/R̌�^�I`��l׺I��4��U��b>G���2ɐ�ZJ��)�s������S����o2��Bܖ�n��~GI{�ʖN4����k��w�5�]  J=G���i���zu/w=ϛ�WXǃ��L����:�uy�2Ch�f�ú��6&��֧��^����ee����2+�xT*	����q����)����W��ުJ�p��,ʼbv��!ńm|ϴZ�9QX��&����h�g�7TK5ͪ�d�f��ߺ� �֦�u�3f���G]4!+��w�f�7g��4� �T�R�|~g#�w?9̢"i�pd1w�N$�I���K/ ��<���#��	\�X�6�.�CA��mH ����k>��S�T"]c�s��#�ѦVn�ݺ���|/�����������9I&U\z$�2Ym��M�K7�B���E:��`�:{�g�lm�!���kUKY:Yz4/�A3(