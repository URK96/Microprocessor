XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ѣ
1��I��ƿ��8��A�ߙ�ُ˜n��91Na��G�s�Ky�����\�vbȦ�����Z���ܩ�Ey>s��$��J_t=��~�4%��9Z�D%X�-g�� 7�%�˔�۴������X�p�a���m�M ���&�8�t�zb7�꼋��Fw~��%��m�*�xq���/d.��W8q�9l��w "hF$^��#��k��Ra:�Đ\��~��[5��Ps/�f��a%!H��4���e`So���|b�ȩJY����;4f��3����}CΔ�#�������#d<�3^/�������ӛ��l��V�0/�BG:{D�KX%�Y�Hl���zG���7�'��Du����Y�r��U��o5��*$��&�M�l� SN���fl�m�!z��τ�s��$���$o�R�_i&|�������u��@�N4��%�����	��Ȫk�N�Ț����@���H����&�Ӆ�}¶%�adP���� �A�Vj��s�E�-�Q8l���'@���S�NI��rU�|n�-�k��P���=At)_�\��Rk�$MW�m��Ĩ��ܻ����{;���ו�E���v��vb9��J�=Ü��sLW=�v�P=9�t�2�Š0����cX%�%��濢��$���C˝X5b����������Y��(�#H�A�5%j��o��/�⽗b��dF#ś���Ѳ��$�?S�Mg�2؍W>s�֩M�E�XlxVHYEB    23f3     910�^�#��.,�±/���v\#����E+�U�$	�hhoN�_�h:-�k� �~��>
g7hѨfbh���D��@�Owy�t����p��9A�W�U�Wi��)e��k��00�k�Xl��I�8����������G��{���f��A��m���b��Hf�M�Wz=��R��h��Q�7E(��Yp��s�{��NO��/�_*<kxt.�F#uM:�}�q-��`�L�=�@�xb��M#P��.-XT�O#qZ�}��˅N���ƯG/Bبv�]�sZ����10� -=��U�~���(���_E^��բ�=ʡj8�����?�C��4��#!s�[���R��Z��=� ��2�}����u���L�h_(r-!��N�ߡ��Mq��W���(S���'Y�[�*9��|c���N�q�ƻT�yH���KF�lV�ӕ��]VWx�����^����+]����7�����ȭqBf�l�U1�2){y�4@ 8\�2޾���G���m:;��g:�Ą)&���m�0����,>^��z~��'�Gq��M=�����7 �(P��
���T����Ҩ��P���1v5�R)�VE���P�����������$`���ܩ���dyvSE��j'�u�J?�j��7b�L���M�N�{���܃��kb�W��d8�`�����L��&=������Y{+��t����U�M�E�i���l�K�i�eG�lu�c�xv�
_n��^����K�ngHaTWإf�{$ltS(�&���c�#�P#�ȋ��:6w��S�p��A1�9)ֈDoBg���%��O����#}\�9��z��X��l�x91]�r���{������z�􊺿6�=��x���~�,�jP'�����Ȯ��)LT� S�#��hC�V�vx��a`��jcb��?F�7���)`���yynoΙhEU�Ab�q�w�YN��?�K�U�s��F�]OV-E�
@������&&u[؜O;���zk�?������)����&�,Qd�ѽ�Ő��w,�
VI=�YQݑs��^�F�.F0�8����Ti�l|�j7Y��~��U1W������h�Fύ��� ���_��ɻ�c�z���N;�;P���ѨB�gas���������g<Z�¾Ǚ@t~w�~3t���mćȜ��J�ڑw頸��8x�`�<�X7������}^�*����ͽd^o(�')pB�`؃˲���VǗ�Hb۟�o%5�P�D���Dy{Y}��]P�Z�9�n�[2E��+�w���o�$'��b��%�%��j�ݚ�}V:��,d���hn��0�(t����Kx������L�"�~b�h8Z�+_pª8�>r�%Sh ��X�A?t���3�����~�u��cS�J���7D$��OG	��<�@!��i(�g#��k��]9)؍�w��#�ǭ/�f ��m���U�i7��̥�tLЏ�.��q`<���R��+�4��!���D�g���묹M�^楏���=�m�������b-+��8 V��!x�R�9	I	����g�yz1jF�4¶�ʲ�ca���cX���-Epc���h �(ҿS��x�ᱸ�G\��"Ӈb�5%�h�ϧ�6�`U+~��2���IL�6�e�V�}Ɗ|�z�5!��O9-��i���Qh��6�фOIU��ę���϶�T�ļR4��e���^���;<'��=�	Ȏ<�zoVԒYF�j}I�6pwH�p�ey�'�)�J.�,�ګe��N��¤x��.�qN�57���I�\0f"���ˇ�%�c�B&!⭗K���:b'��)@�P|�c�xŤC��$]-��� U���L]v��qGo nW�h��	LՂ�:�V�¬X9w�ۖ��q�I?�n���.ÿم�V*dƅLqWmJL��1��epQ��&-k�(��~R����=2��N�匑���/=�	���!q�͟���A� )L����=�;#���I���y��1��b�Q{}��	|����!�1L�Dj��Y�����E��o�#�M���;^go�� |��� ����s� ��~��Ć8.�E�[���9��A9���\�`�(��uo�V����;?@��84U��zU�1B�7�0|j��I5�r#�FKzv��9߈���k8����w�I�s�8���2IC\���Ǡ��'-��ӌ(%�\U�5��}���P� �X�*��Cg;~��f K��]KtOeg�"Gº����*R�:�v��