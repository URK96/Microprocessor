XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Y�I��F d:WЃV��a�+CGWzc�P��J9�Ԗ	�$xC����1��5̇"v0)����A(Kd�L��&�v�l �?���k�uޑug��xձPP0_-�pc+ԅs��b�M)� Ȫ�P��|ǖ��R��	��V>wt�*����9GC����.;g"�)��A>��������v�֎����� U��nw:�zn!"�e M�`k��:г�_<s�(��d��=B��ݝ���_ ���-7g�2X�0�V�^�>x��|���5[�Ifdo���iE�Z3L�U�����ڿƙ
� "��RYx���#��i��p-Nu��u ÷�	�?�?lB���� �� =h����q�="��h��L} @���}R,*��xW�Mf*���z0T�h�|���_�����]�����t��+w~�����D^�i,XK�c�ޝ�@|xk�4>��G�����D]-z�P6�2܈�˰
���ZΛ�\[}���,�>8<h����8�.��E�w�P`H���l����'�}�!jq[�t�0���o�{����7sp�*�J��u�wo����+�H�<�*�̨n���+����7�=:�S��]2�>U��f�7v���b\�U`�zJ��ɽ��F]B즿"cEV�K�-1vp�[���w8a��H ��ܼ����&o��)`�A^� w�����Y��Ueִ�.n����t�Cp�nRu�
�:�l�*�vݦڰŠ|�i�Tn��y�D�Hml���!MTF$��l�l��XlxVHYEB    d88b    1610�b��ڐx��~�E�k�N�����텅K�e=
��{��T��q؟np
|f��b�z&L���nl�j����v��J�E�s}�k����Ym9��{��v��_�y��;�svq�j���s�2��)F�,�����7�5�8<iB��u
C�9���m�HX�]��P�(6����>�� �IU��@�8;s�25x��_��m���Z�W���ttwr>_ӣ(G%T3�pGSm������Zgπ�{c�Nj�p�öq�[�� pA���N�s��w�&c7���c�گϴÜ�8F&�;¯�݊&������b���^���`��r�h}�"흕�^}�8c���dG�J/��>9m���0�����0�-��l\ڑ��,���^��b�L�<�_��,��X�L��5�aū���V����M��Wf�A������J�k��<� ���`�nԝ(n�D�����qǝ��\d�'�:��{ *�z$��Fu���X��+	d�(�}D9�D(�6�*+゚�u�0�h�����$��w�n�t�[��l������н����8�gߎ	�>�o���W��P�C@�TX#m)i/M'�!��\�$X.T � � ���n���l-�ue����ӗ��S��"��RT�r��N��I'֔�2odL��j�HLn�"-���I�r��#礫YMJ���=h݌ޥDn�}1����>���d�q׈0X��ޕ����n�������-I���HA�,#H��@zIhD�Ք�#f�P�)�9�r���>3V����:;bi͇��f׼B8���(�{ø����Y,��S�Cޢ���lv�1�;?�|��-2�e��3��n�>*�ߚ�,��<���2hZ0[H`�69"�3Csy�\{x� ��!�e%��B1O5L{��^���r�P�տ�w=b> ]�ٰ%��XFC�n��@�X�A��>�=
�a�I*_��H1��wd��N��,4j/9�yuRD���-���@�o�������/k��.m����|�8@HZ'�� �-��TU�V�u��*No8����'���U�;�q�� |�;���X���IqC��(� �)��4���ToA��p���
�o�!(�=6�������9�n?�8�dUs�,���s�OYŚw���f�aŝ��z�,�!e
cVMxG���:��	�:�	7���A ���3\��cF���#�`h��q�wf�/l>�r�ME���3�Bh���>=!v�[J�&�[�DT/rX�C�xX�8��yf��۬}o�[��0C�7��l�"V��ί��z�E5����
�W JИySu��>�[��xoLq�[
���V��(H_�L��7+�Fh_w���
���ƥ��~C�pAھ���2��2�Vė�i^����]��F16�8T��6 ����G�~*��Xr��S�l�%�]�'T�ϧ��-�k��|�^{��z�Ÿ��I�Ф�nV���sm���{"�S���Ү�V�oC.��i5�S���z�C��$�ӗ�S����4��,�j�J6�nR�f�8���X'��<n.�^�NFS�'�Ə���Hj�;��H\��a�6�`�ǈ�������:D�"T�>��K������~�>�/���2���h�Vh�ΧܤU��L}ˉ#��|.}΄RQ�DP���0M�����#~-_�[� ��v��iN���o��ḏu�ܽ��PzjK�:��Q&R���z��!����Fh�Q#,�\��G'F�$X��_=�_ �� e4�]�
���E�dso����=�Tʑ}�������ю�̺C�{\�u�^�1ON���c�����0P�$3�t�G���4�?�U�ou�r"��ܶ�A�=�]�x�"�r%���U�Z���;[P�o�(Q�(aJ��ٚm�,Mn꽿�w�P ��W2c��d����uʏ��B�?��!�I��Cv筐f�|3���Nj�JۖDԫ�䋵���ՙ6Z���))e�G�Cf�l���y����6@)�=|�tgStCmi��p� ���!:iһ�3G�q�t��2�_�J]f�X^�@�����i�V�H*�j[��A����q��l��H>Eii��3�R���'>@r\/`a�C8�S�|N��L�Af0R����|�&�bY��4J
Cj��g;H�"�s��f��=ݘ�;?�3��/��C�'Z��E���:gs�G�r����`�[��m�0I��t@� ;�n�����w�>,Yw?��>T�L�nb�z��P��=p%�X̎L�M�˲|�WX��l0�p�.hw��P$����e;+��r�����T�m�������jyaC7������hQ��6����iT�gu�+M������m\<ӡ��Dp�%g�Ap�+@�Kd���%�p�w[�8�B�t�����٘v_��n��d#�\\�Lu��t/�r�AKg��B �3Nlt��-���p;1��G�,[�_p�a�_O#���W��Z���pP����s՝��_��)�)LI^xWa3���/#nIa1�A"����i˗��{���&J���6�;͂'��G� ��m:�F
lT^s�0��k���Y�����D�=/	;U2�W8��o`x]D��k���-�4�`�]v�����;�������l��/���Ҹ���� �%��� dBFuq�c��Q�l��������
]����f��F@a�]>$u��޾9����D���5h�EC�$2H<����s-3[v���v��p����eBܞ��o0L8�[���;:��m��:]���ƒ����=h1��Ue��7E�c�D�$d;Ԍ��A
#E�p�B-�_F ���ٔ:Ңu��M��6q䛝��r�������t�2>+s[@�%�q�x[Q�O�C ���ahA/DN&�^�V�`C�	��߯�-��3�j�/�p�tm(^�49�P�B�����(g��~$�z�9ɲW���7�p��?)���-�]��,��s�Ck�>�\^�"h哯e<1pr�ֲ���X�����o�=�ɒ�)��r��Ůk4���7#w�^��p��m��@��>!]T�9���N�VX�Yۘ�y�����01�䣙�2�����S�F�؂ı��?%oԃ������".�|yDw7��]���3Pе0�~�HI���t̘?�����nb�z�iDiS��X��
z�pn�[i���딽 ��vz�f/b���i�R���U~H�Àl������{��f���ՅE���:��0z]��Y��`
��R@�g�2��E<��Q�s�x4�rE~����E�<녏�]ԡJ�C۴'�(vA��hC�yzo�\���=���n�Ko��v���!��,�y�k]���E{1E�f�'pq�t�~!#�ч�K{�-������y��~E|����)�@E�tE3�6j�i^̲��Y�d��򔂥/��+�G$.�|����X�j�򔌣�''8U���:v�-��òy�����Fg�6>�������^	�Q�U[ɗ�@�ZQQ�*�hM���G �ee��n!���j��3��E���L��3��˳ʣ>�/�orP8�)/s5�
���sQ?e��i4te_��*r�Tw�nJ`lIj��(�Pnp�]Ǯ�� i>t_,e	?.���([���.bz�}�<�������(���5A;���&f(�^�3�9gZ�f,��c7���ԇ!�F�ٕb1+�47��<����B��`[|J��P#%�(�|kSr�����;JF� y5σ��5stF�y�K ��ճ�|�ؓ��S:�J.��7L��� E�U����,y������~�..�^H/I}gIRp	�s���'CI��-��h�ϑ%��LעT'��:'fO�c��jn���g�;�``�!�7��x��ܙ����qu��V��[��[�}�m����M+�2�m�m�Ei%z(�	���E���S$8S�D��������X����H�-r<�����
������k��E-���"�LB��3x��X]߯GS#f,h�*�/��c��{�JJ9}Q�N�ё4hO�H)4}�xa�G����ƺ�&9��*��Ox ^������] J�F���L�R�P)�I*�^�ϧ�����	���T�����cUC�|;+~ ~�Ҹ@�ٍOF4f�nP?p��t��r3kzvл���@�>K<�vF����C�c���Q?�Fg4C$��7�+�A^�o+�o�r�ϩ �
���W|��;jM�ԡm�ǇC!���En�eI���z��&�%��@=���3�����R���'B��3*ɼ�s��E�68���h��[�L�x��c��_�l+S���i@�ZG��t?�t�L��vӯ��@�H��Y/�Q��s	Iٶ�YH�osC!��⸾�u1����4�����,)/���}�C��	e4�w{�0P��l�ϫщydNrF%F䯂�Ka')��A�e�O(�ύ��50s@�����
"���cjob�:^+RR��"-�c�dÑ��W&ڐa����*�2��z��I�~m����`���?�Ն�*�<����\��}Qu�4��ú��M��,Թ�=�T������»�-e�<��7=G�S �ׇ�7������7(�&-�'�E8��b���쬯�:*���Ӗ���#z�����).~�r�љ�0��Rk��n�@_'0�~�(���t��C�ZkւBi:r�o��(Ih�,���x�B7��qɠ�K9:n��G���s���פj�	o �*Jv���)�>��_=S��35m�J:w���[��I,�:n�(w��\9U/njMh,v叓�P�Z7�^��I��_�y�,�{�z��bں�:�ͷ��K�~vD�YDT�|q*�*�X�L�8O��^��WF!]C���K�K�ȿ�Z��gF^9�t�m�����Y3�;I�-�P�i��,���@�!�X,�(�Z�Őc^�W��T~�y-U�CQ��eA����\�6NW�$*���n�C��ג	&���4�Gc`���D�D��X䟱��U��>�~�(�t�N��`N���o��V/�Ž��A���iu}al<�@���T�a��  A�Xg�tɟ�:��vS�J�4	��SO\�'w�z��DK�Ӈ+]o����Y��f�Wr9�\6����s=P��0���^?{N0L��Aaaa�^�	�����Iݾ��빽�5�Ә?�K���ay����7_7��3��Y O�ޔ�Y�6��Ѣ�P�2<����blU���q� 7"ON-�g[d��u{�o�q*P��;���S��r�U�#s�.@٠��Ɯ����NdB�t+���* �Bw�]4�-���y+���O����ӝY�;1/O��<�2���`�0z<E�C;����b�}�[�:CD��٦K�/$�UQ4�<��B	
n'6�1�[�Ņ�]�Vq �R��*Η���x A�FN�ח�.i�{^~�lČR���v��0DGH_/��Js�)��'�/1PaBB�ܧ��}/�i��