XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���3�6e�ዘ�6|���L,
x���	����yj�8�O1��7岚��tjąwK];�A���K��0H��Z��AOT����K��b�������+O$t
Z`��$�6a)>�G9�X}Q���n���t�x��W#� t��3�K@\��̰>R���C��p�hˍc��T˗�輰�J�PZ%$�Yk�eQ���CRV�j�� �����¦wT&���8ij��Q~�U�:�!��/��d)?��-�to++�g���Cc�\��]�����Vd<D�O-��O��>��Vc�Nn�����t]��[�U�p�1f_`��'�\T�b�9�ݗ���o���׃s_�р�R�j��W�*����;A�� ��b	��l?�ڀV��}��U��4}���վ�,C�����(kF\l����쳜}B�(: ������ͩn�&� p���ʝ*W��[r���:�9!)�8�������wL�_���eΟ��lG	�-=j�tQ����N蹒��a�(�T��*(��o�Q>��7һ�K���>��uٴ/!�W�����L:^�kq0�\���1�T�]9��l�g&U�S,��b����f��Tѫ,�"ΝWde ���&u4Pۉ�7g����;�Bw)����ķ}i�O�ͺۤ�Ϧ/U���7������8^r`1�2]E����_:w
�h�q����3=�V�́�X�nn�J�Z�`�����?�qq�C4"��|W��vi��f�3�-����%G�9\D�!ݹ�XlxVHYEB    6408     e20^���ǽp�h_M.c�-?�|�X��%��$ 8��T,��	��k��В�*:��@��w:���Ȥ�p}lhk�`T|{"�)�f�����.'�Cfm�k��#��b�`v<��3�ٞ�wńl$�]e��F��U%l۽�E���,F�pvG���%�|�0�&v�H��)jP�/~��=�֗��DA�Y�LI C`�7c��f������1Ly�e�Bc���D�P�cz��H���ϾH�UUV3ٲ7A����~Ng�u�
UgLG������z��6x :i���* ���x�̓fo�CA��o�	��YdI��-�9���=���4���e��2/�h��L��&�@�p�V�ǀ���������}w�J��z�2�Zj�#��CՆb�YT)������Rm�n�)�T��[((��RɊxEG�X(�����&+I >�C�zf�����Yy����.����`.s?���J�ƼiGzw¿a����_�mc>��>�IgƖ7\����S��D`����]Xn�DT΀�H��R�h����|�ļ(λNǮn'm���0���a4���%�S�[��%��bn�![�x�
DF-g�Z\�g�(��4({�N�3%�,[�O�u�!� �"ͪl	�xҥ`��ֆ�cGO#a�JUK�
;�$�^�Y��n���]P�n�;^2	�/���l��!MTv6~b�%���-˫�����)v�]%�ܓ�; ��z��0ɞ�$� &���4���eÙ�t�-��@�/,�uB�j��n��<�J��O5�<+�+{��"��:X׶k�d����_�T�)ө1N�R����̽Qr�M8i��t0άRn-<3.i¡�B%�"y�ͧ��\�RSDT�́<�pǕ�>��,�����T�-��>��qCm^������bŃ�9[,�^�s��*È�-ԁ����/�"��ػ���� <�n/7��'-��
:ť�`e��=<G:Q����	��=��} yI4��D?'V�x���'���}n�JmJ�Z]�㜠�'�\6�b���zm�L,kRڵm$S�ż9�"�$L��s���A)�F\kxz~��q��-F��d���Dߎ!�Sy��Xq�7�`�h�nqu���S,<��[,r-&�!l�y������T�����U*H�ی[ � &�����H����֯�NhT��>6��c�1w���g=`�`�ظlh9R�o����u~/�z�N屇$����P)���%xpuN6�S�S��Y�&t)k�N���>q�}x����6;m��}I3��I�в����V	��;&Ά�s�t�_���>_ ��)��y/�{��[�'Y���+!�3�;�%^17�@�z�ƋvK��6�[�80Ɵ���%� ISȎ`�ю�9�ki��W��2��o�PV�d�_-<e��󔁻h� �?I�����E��)��&�y2�4�bu�=��S�k(/Y��H0=b�+����~���ih�dB��m��4�K�W`V[�,葍���q�g�^J�`��>�y��fo���
$KO�����*'�y�8ÍTbb ����a�̵�Z��-���ݷ�}�!��W�T���V���9�x�~Hq�	7d�"��o����.��^�(�I/HH��P�f�;Vӵ�b���9ȝ��f��4������j��`R��z"3j���)�ƛ��j,ZxՈ+�,]�.�,�"{�2Qg?O����Ӊ�a��n��G�}��S��E�=�<�L���8��0�
.��7^2�#k�TM:M@��lL,�ki��]}��{���W��Ӳ�[Z��F�̹M�I"&��'��r��^_\��&�����{�͙E(?�*�Y���0Y�y	��
"u��:f��FeT��s��6A�[�����?t��k��9����f_�u%o�4��[�V�ƥGц�����~J_�'�L�lVF]?_��m&*��h�x�	E�	2��R�]���n�/a���{D�BV�PA#g�BzxV.tYSfTo?�4��������Bʪ�K�P,h��A�t��v�����l�#�!�D^�p���n��L�˅JRH����#�J�� a:�쵿�l���z_�%����5u���e���A�1L�L'��������K�[��O�t�Qg^\�r���uq�����}���?y��}���7Q��$hN��|m���2�Q�7��.�w�HN�O�������okt���J��ⱒ�53Lm3"�=��|�^P.,h�gՂ{��"�S9/�)J�Ug�wgV5�{�#�(��~�:[2{K��u�!̀���o�ł�8֍(�`�W<W�^����񅆺���q��C�-v�D��썴��fz�	�D��J��c_�u�\V�V�j�dp&��`�a���&L��t�Xbψ#4U��.�g24�\��g	os��I[�&�n~���������e7$31�^��W	$'���\�I��Z�+�e!��g�������\�n㒙²��~�"A�{�ȅT�N��QUx0�b8��,$u��P����fUY�'�5�����c�7&�b?۠��b��*7,Wj�I7}D�@6+a׏��ܗ|��d+�_�L��8�ޘ���ź;�O.��F�k8��*9/�0&d�
�t_�m0B������� .}��9ʔ�o=�1�Q�v�[E��W�z�����vi�������֙215T���d#��f���h�"RE*c�鰁��P�c�7�U,B�#�A�ό���BM�nl�� j8d��m��zŇ��i��8m;Д�v֯8PƘ��|'\�W��j|�t��nηV�If��\�W�[�cDwT� SY�?��4��}�� QO׉맴dC��|{�
��25��Jh	O)�-��⧂�-hC^M`�p�ht�N�\x_P�':��/�孹��s�K�2�	�'o�%/�T��]�/�Xm�h%�h�F�Uiˡ�k���]yѐX����k�{{�Y+*�n�������ʽ����I�dD�l�~Bן���9��=|&�ʺ��_�$�֦݊=�5�6䚕��v���9��SN���*�hY�ੇ��k+G�eT�q�"{����e�my�/ü'�~�!��,��AA+%�"��y�[�Y:��+��&X��LoCL)R D�I;�,uK;B��u��:Q/�O��v��6ɩg֫�pGD
rƵè��t�
WiJ�9�%�ی�Y@4'���M��a�t)}x�����J��SԷ�zf�e��>�N�3:�S�	���m�ru�`�5.����&�U���}Q��B�O]��L;��}��a���%_�g�9e�a+���fDa�v�mm�`����u
�K��Ⱥp��ݪ��)Y�l&�cd�Sv����״l�F���=5�WJz)����jV��ydK^�� ���2���%I)�C����`�,֔���捼��4w��T^�ȅ��� ��98&+�I�B��LE��
����#�12ȳ�����wl�>�g��� �Z�H�Ir�;��8M}���qo ��^#ZT��:��O�b�?�G���9C�6�[U�[�