XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��AJ$�<����_P9��[%ޚt�h)R)��j��x�����w�K����B!>'�]���g{L��,��H����<�I��Q�����ӧ�6�d�R�,��s��@�Sw	���~u�9�J�F���:���n(�w��]~m巑��� y�;�Ҁ� B�NY�@Ђ��N!֔4-��]�����6�0X�
$f&��JGv��Q�4ޛ���qޑ�O���}j\.�[��vÓ%��I<�Gb:��w��:�sa�B�b�xd沯��Mw�#XR�:��(��V���1̏��|}
 k0�!�Лp�:kJ��K����6mi��a��#wjYa�bg%���
�zF�Ν:�и�pz&��n����F��>�t �aE��{����>��=����X�=��'Zf�m�Y^�0���᝞^.��-2�j���d~g+�dG��T=��;����3ы/�1�7Ï��	��~4u]��0h`ibՖ稳�ͰZ��<_�1;���i�p��c��6Ț�f{u�.i�]`��wݒ@^[#g�CO��a����w�D�Yn�l��u(��9��fT8�?*�j��G�:#]�2�7` �5��$N�#��$��/�����b��@���{�$ڲ޸�)��y��%h��`q$�I���?䅍�D+��<�@A
�4�����;�
�[�k����ڶY �h�K��q�;ñ�����RJ�:�5�1c�@�HZ��! t0��Y��O"��~t:�g�,rXlxVHYEB    26e0     820��*��:�Z�������1q��r�݅�EC�Tۗ���諬�ZP��Jh4'D��Y�^Q��i�>ҕ�0��2��g��������U@��X���1�|��BoY �78�Xo�3 V=r�@q	�2��ɰf�T��-s��"��B!rlѮ�zaB�c�w%��Bs�y[RCr�kc��b��ʺ�`�)^�8�p)Cn�ኗt�kkyBZ��?i?�hvV��"E�C@sn���V@&�OaV�Q�%�z��I��\+�7I	��޶E�6,�cz�r�;�?���@��5O�ՙQ�U�w`��F&����1h� dh�x^�[`��'�&�A����]��&�Y����M��i))�8�+r:V-*O��"�#�M�?L�����&LD��n�Uׁ�>��_k�͑�|��l30	EM����>J˳g���n6������M�~����44ö�;�o�Q��6�x�� e����T(	ב�_��� k��^Qjg�i2�Pn;�Z�ډ��v9dhD<9�f�ë߭�7N�>�?���q�͎a7˦oj*R�1�8��Ê������TC2�Ǿ'[��]Լڱ�����m	��_5G%vN��*v��3��2 �J��^�ld̒�����Yw�B�<�q�&M�^�*���X���b�"���
zՑ=���h�ՠ )'i�h����0FB ��PV;fE���V�O��Z]��kEHB��>S.1���7��A_E��oi��=���Q�� u���r�qF���!��ў��Mݣ){ρ���I�X��
!��u ��26c@�%$BC0E�(N5�KH���m�h�m�r�����
i��Gg<݄<o(V4��\��g4k������P��a��o�Gڥ�%m�[��Y�2��(Y�H�NB������R\�~��j��8;Zm���%��!�d9Ek�&�c��)E\#"И�'��Z�i��3P۩�:�;Ƀ���?b	현X�Q���_���:���.�w7=�=����t'�9��L{!܈6�@{~�  ��U�)���ԝ�>����9���΀u��J��2�;d�QG�
P ��
�%H���-��êi%S�^6����.H}{�=���85�@-��Ds��IJ������X��L`� EW'(��d� y0��yl�7�xq�����V��O����婾����P'7>��g����O|��ڊ�yYMǄ1�s��Ŭ��>
n�6$rE�5��诵�Lw��ʢ���N��^��%�!!�\8*��k_�gt hn�ҕ���[�Ol+��V���0>�j��9w�yRy_�7#kC*#a* �o�ꁙjZt���?(�W�I��3�A��N5�m���|0æ-�fI�P{m�#Y�RS+؛fw�w:��f�g4�+#�H��R�F�C�6���qz�x�����_�,o���T41`/��4E#?L���=��Ǎ4
��_������V(BN���9��5�{�9*"f	7�4y�+�����[w7q�}��ť�_<{`��g�)�$G�8<�Yx W�Ӵ$��[��*�π�3���(0K&�h��Z�;�{��P-r�-��oj�&��x%��bF��}���Ĕ��Q/��D�l2!��݄������s�@I|��Ru�mb�g6ֱ�)���L��o�e/�pG����m��k~�Mz<X��eZ:���RΥ0E�+Nn��फ़�y������!�=U@�o�~�5��h�W
�N�a��(�c���va6�,t�&3y+۰� t��xN���\�d���߅^&Z���0 B�	"(��M�bl�{;���ƻJFRݠ4�����Q�̾t��X
�+M�Q��:�xv@��_�Qq�����6��d`�|�w%��x�����5����9���h��[z=���ϳEZ�cz8��
�C�)�:}�������r���X�1$���!?Wzv������;����x�ڈI7oL�~�7e�?Y�"�� $�S�X�?���2U���ۡ�h8�?g��Q�ǘmŝS�P���$I9���46�O��L"�W�L}��