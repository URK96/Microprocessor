XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Tn��V�֊�\%�
�6�P����2�S��*t�W?��X��.!����BEdP�b�@���{��p����F�v<�Z���\P�ez�D���(���gG (n;F6�����<W�m1�������$���8�_Z�K������
if��D�`�������]K�2��$9��"�/%X�Lj[u�9��z���0��"n�(\֠=;�=cDnq�%��<�V��@���0��Y��,`R����1��8����5@=�!Q���8�X0��6o�R!0(��6��ӊ�#���}��G��TwR��2�}"��j�P)��w�1p�H|����>{ [��gF4�#�6v��FG8�@(�>�1!<�R@�9��'䬨�P��5��z���Ow��2@�T׷��9 ��:����T�:n�R��c�E���)���UW��j���l3��v���!#��J�f̣�;LbĘ-W\B����>S���(��&�Ȩ�W��1�#^/X~��c��"��t�K���"��F����P2N��m$�:"4<`;m���f��x.-�I���9���(^�^��/ɛS%4�*˒�k�v���J��dOvk�;@�L���娊.h�� X���n����f=���l�]%f�-����'@��E@;٠���H�@�Zaws?q''�'�䗟�=�o� ������M,��7�,9�]
��%�4�AF�Q�!��X,Kj\/�ī����4��h�dg����g-8Ӛ����~�XlxVHYEB    3a19     d40ߺ�.�b(	����]C�>]����:��}���{�䋕nNCa���K�E2��z^�^�]�-+;?7`)��h⬠���YU��-�M����L����q6��`�D�so�*�R�]iw�q�1�BdpW�ڞ���u4���7W�-�@C+����� ���t!]��E�č�?�-��n��$eM@v��~���
��
 D��+� �Z��B$��kv�2�r��ŕ�.>�����=��E��p3�B���\��a��lS��U"���0 f�C���Y����� �igW�]O�� +�g��J<I]���h[RA��1��M��3.��B������ �Vo�K��(s����ek�U�M��Q��{�b��f�V���O-�����3:"�<O��Qӣ���i-̤���F"3��,�Sv�Z'I[���̤_���{�Hk}R;��]��hy��R��,PF6����-�ls5� �w+����&+|�Ģ�{.T�ϼpV��hw�o�S2����zv�}�'�¼�����ݙ�P���M��~.�ơ
N�G���h���@_�}jC<,�u�����z�x�w�nK� 1��0���փ%��h��aSa]�R���3�t��5)B����|��O�M
���q�wn�F&�����'�0���7a\�!�J���qx�i�D��.�.j�.�esS��߼�����E�P�Ի�e�;RW��w����(��;\���.D����I3�aL�YL�;Y�֝�4gpZ-�ದr����ݫ��G��J��/��4��X>k��O��F���Q�@A�p��Wp��<1`r�)���f���T������ve�#�3�*��_/��|a�F����}��M�{�����H?<�CPp���<����C�1�)�r��z߇�i�dV�Y�y����)B螦��i���=��{�f,˲�V̥`�l%��֭t�g)>ۘۘ.2yK�.�HW��5� h"�yFhy�B������X��j��|g'̌7r�{�ɘ%�:�|Z�=�u(��&�Ɩ�n�&PBrt��d��b�u�
�6�뾽T�r� ,��5:M���n'}۫*�
q��OU
�`C�V����]Z�ۥz�c�!:s�͑��6��XPp����~��d+�D�U����_�@�t=ZO�sj���L��ͳ��|�Ď]�5�T��qp����o���&�4�T��P�7���Q�g����͡��|tB�#�7/�5�j�>�s��?o��]��} -�������Z}����Ԁ/0E��e�l�&����ǃ�����=ٶR9le�vY�x���7{�����q9����~z�F�^PL�k�'7N{≮�&�TH��/�K��eL����7�E J�/�wZ��9/?��d���/�\�,�E��$���,"��Ϧ7������s�X�s�&�[�1B����������FRTs���D��Gha�}��U�s���1	k
o�a0B(���
O֙Uzh��� v�;��Z��'��T�Ε��'-i׻�~�'9TI?4\`Nd��4��	l�x�ɂ �/�]���[��C׆��Ƙ��Q�X�A�-@k�m�� p�3�-���R�����9���2^�>OO䟹Q�eJ�f�¸c��큼��5�~ٖ!G�F7P��wt���9��|y�T� �� ֞��	���"/A�ҿF0m�4���'��}���'�<�x���i��6�Gala(���r�H}�W�h@���Dh!ѨJ���!���D;DK?�Yi���ϩ�2S���<��i�N'ܖU�?��3����J�U��l"Z�i��G�Fݤ�(s�7�� ��W�b�*�w�b�eH|q�-j�jmg�l@�lщ�ֶ�m� k$�0ܙv��x��I�W{Uv�r��B��=纒���R�P9�tZ�5���^�]������@b��#�x�@��Q�C*�����pȋ_:wIoP�������e!�O��x
�5?a�0dw��lvuȏ�q��W��[8w�Ha�J/�MC�%q������O	�;����h4�?\�R]����:��
չz7D�B�{F�����m�ȋ'���M -��(�v�FJ��iW1�x�rR@���\%������E�z�{������dI亲۟72
��t2*�n�wڃ�%�_V$x��j���:#@��]İ�����}�H�UZ���w$/�(�k���bC�yHNϦ`r~Hb�Q��!44�%��Ӱ}5�V`b?U��W��s��]eHM@%W�g�J/�!�ڡ�٣ C�۸����X[�}��+��Æ�y��J1�}V_�K���R�3wSX}>'a=�ɑ0��y
mql� ����Ļb���|�U�2rGP�hu
Ͽ�&at�K��|������6�Fp�2e`�F�_xo����֚�u�g��?���-�\���)�p�S��i�x�!�3��G��^H�{]�����Z 8����	@�Rg;�Y�3g��b��I^er���Jl$ �2ҍ$a7�3]D��`���,!�F����m������l��e��MfF�p��$Gp����p�>�V��Lw�1��\�k�oɀ��ąq1��)P�3���a�B,��`]q���*<!�87ܴ���Bu��0&�:]�5���m3�>�p����!SQ0�(lECZF�s<�����/t̜�絠}�\�E�+� {�ml��^	�眺6�f�.K�,dt�T��۳�j� ��|?��.�A�e��G F��)q.����Ѳ���1B��j����u�n�k �ߟ]��V;��f!`N�k4��h�?h8�yc&㼿�	#�!�1u�)��v�qz��N�M��ڻ���wp�F�A[/1����m؂P����wz��߸h�J�2v�8*#����Ki�|#�ȍ������#D��/*C�0�l�5I�+}�|��]�6|��#s�_ƾ7���ܢ����F,���1��#��r˫_Q�m�܏moQ�L�e���d�ա�;�7�v׻�̇;��m:�Q�`y�}TOq� Q�.�=�����Q�����7;G����
���6�����9��~����.����e7$*���9}Dc�Sػ��f�����[~�_Q��xJ�-\�\���+��N	ɰT�L��R�=���dE.��Rv��C�,�k�:��S6q�A$%�+ H��:��@��J�9N�P�tQ$���/k�0���^U�ř�(���*��g���v�T5`ƚ �����T���o6t�tN��Pi1��B��Udգ�)���37Io~	��߭*�kH���j�7�U�����_"2����x/m�$g��