XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z��Z��PY'fg]�.����{����&;2f�w-�˽aW�>��X����%�z�1Y�͊w�.��ĳ�G�fb�R\�v���h�r��*L�Z��)g[R���v�[�"�.��`���"�(�|Veө�Lmg��p�5�Tދe����E��� 0�f|B��#αz�1���&�b�$X�Ve�I��Qz�JHI��*,���&H�y��(�]�yf?��d	��x$���}!Q'{�� ��*��`��7�?#��tZ��`��';<c0L,��-r�.�YF���WO]6|��ڲ�J�[�a!n�b17�׉���C8x��=�� �	�%�_�J�������֕�3Dެ��]ܨw�Q���֠�^-ZR+��jz=+P������u��9�8���ϣ����
r�'j�.GN�i�A�/�M���������"�]���i�b 3X���*���I*2�X�H%��I��+ϴآt��h��mXz^���\�T�5�u x���9�a����|o�A��B��b���k,jT#;O��᥎qB�������=.� Mv=t:&��-�� (vm�dV��I��*�QadG�b+8���a�q���J�F�aUEiSC�F��f�18�#�6�zz�&B�@3aJ�����8�G�_/B��E�iä�GO������p�*'�'.W�=q�{�l�H`����9i�$Y)X��Cb�^Ro��cb'�z��k}��Z�j���$:����*�e$`2d�Z�XlxVHYEB    2864     8d0�y���Ή�������s�¸����rj�ޱ��+e1��kKu�DԿ�m��.����|�H(�Џt��ȳDX��R=yiC���	~p񦎅����}�����u{�,�O_M���!�;'���G���9���IN��Wܵ|ҏ�A��tת�m_��OM� ݛ<��4R��#���Y,A���;��ֲ�nR*�F_5�G�^��3M����ٵF��F�gO�X�R��:o'�������D�0�D��QV��'�[ᙑ	k����I� �����č�FJ�4��`)�;x^�n��o5�-��UK�m���Y�����xj�\��!Ñ�ȅ��:�Q�^�Z��+���}W�����ީ�[��0�~Ƨ��pb KD1�w�)����0hyۖ�/�j�i:
+0���0�&��� [�e������Í�[Mo�
�!�.���L���_�@g�Km#���J��<8�		��%���	ܨ�<ڀ�Rޜ�T��.��
Ccf�"���׸�q����\6=��I�nb�m����~b�n)}�AM�Z�L��O��?�)mD�?]�z�E�;�=4�1�������y�]��J�L��x���UCn��W�h9��B��u�=]Z�E��T|>��y<4f��Ա,W��e����;!y��d�E�Yk�E���χ"���y�	"�I���-^��ږ�=8����[�w�N��ߒ��zt�f=�6�)���>��Bx�F�IK`o�+H���l������t	Uٮ-ɂ�v�:}3Ȁ6ǈӅgiР��[zWZn7`���J\,�x���=o���8>;�������}��m���Ĕ���U�!�E���0��M���2a��rV-L�u�,��N}O����c�S�Hܥ�P�v���Ѧl���K�ӄ�DǱ&����ƥ��(s� Ȣ��
4$Ln�lme�U�&�@���{�R~HJ�"��<t�Y�K5=�,���>Ȱ]����|�h,���>D�����tk���I����TG�W;ϥ�t�~ 5֠���B*��v5�q���l;���`3��	sZ<�$	���W�3dp�J~:V8o�$���l�H�t$V;�����=�PhB3�6����X���;�~3�_m��:���12P���$�@�@k��"�h-�Dm��Ҹё~:?R �v��퀝��Y����!K��Epƨ��]MT�k�X���� �<�����u�B���j�D�)Zb�}�3A��\�,K!ڐ�xağG������A��n��(c�g�Vt�K��+��{�@pn�{r���x�-񆰴�%�\4�.�UO|/���f� ���;c�K�jF�h����4�p*ҸmZ>U�v6�ΜX��\X��ǃ9��Df�Y�g�#0��e/��-��v�<ܑ�35�!|��m�lq�cx���Lw��$��zO�.������� 0^*����
�y�:"���:Y&�	�_��� :�Qt"+��N���L����0�Y-W>���7�R����S9s�ړ=K�&4*�!1ޒϯs/�_y �	�T~�{�58��N�T�S]��!���m�n�Y^6�G�����a1�
t��:5!�o!u��r�c�[��&��|��������ν������x�v�Q�q!(7F#^�,+��	j�v&���i�e�!ݥ;�o\T��T�dSGL�'����+�)��&(��JpP�5a�n�nځ<V3�&RaŒs��02��3��)s��p�þ^4��Ga��mj�æ��rso�:���W+&�� ���v� ��W/=
����:qJ=7vB���3�~~���v�������3�QeA+(N�4��{��Xq(�Pp��v,������t��^�#�1�E �6��G�T��@�2��7ŏ,M�Ny6�[ǣ)������uՒ��o� 0�q�h8�q �;5�k党J$�0�W�br���$u3JK�Z���@F�o;�����E�v���x�@�a7��\F�̠H�-��y�x5��R���\\�w�h�5�Ȓ&<h�A�EY�(� oˮ3Q����p��!����l1ʊ��i�i�v ���(&I��������w�PQ��|b��4�}��ë'����Z��N���nd+�Ah��c�w����0¯�p�sk����BF�!PO||ju@�m�H �����66u�������"=���p���=�7!