XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r�à��3����GU�t{p��G��\�#�+ ��jo����Vλٷ8�å�^vZ͔�<�����O��p�E����ę�%7��8� ���/y��R�P�&;{c#1:�� %���_�i���E*�!.���o�zS�c^,Z�O;Hc���E�i�&���e�U+�oe�[�ʯ��W�P������3�6�ig,��M��^p�a�6��9��v�L����0�b��X�[�M�	���=�6o���̥������H��θa����*r�BC��<s<������ʈL��%���AŃ�H�d�V���#n�N�ɿ�B�Q�kU���y��>-�`[z
��|4piH	�MG��ײJT�����Z"W�WϸU�-1v��GE�5m�@1\�y�j���-s=�wd4Q�4A$>�E�Q���m.|�^�-������¯���e��,w�i
I�O�ˌz.^X$FR�R���6�w��r�w%��Z�萐�a�pb9Q�;�Ak��p��-�J��r ��$ta��Evz	�a���e|~n���K͑0������b8*`�A��ȣd�8O��H�=aO:`�')j����5�{��/�W:,�����!cof:������x�9�-�PG��: �3�1�\Lb��VE\zA�U���L��u0u�67���)����?��5a�
Hu����M�0;��G�!%��F��s�'�޾��~ߥ�N⿣�e�K��/�i8p࡬k7��A�/�6)1�RXlxVHYEB    6fd8     c30�f���iY�l
����:�?~��,C�fG�D�~���K��r��/������l�$̝����5KKTA,���u�{��mfI��\R�ہ�O��4�cp�l�_͋v�f�}�Je���*�.�~�řx
��=_����ʊ��*�� λ	�� �8�*B����{�y6��i10�5��u�g�� �����~J�)n����(���-�ʯ8�|j#]�MDu�����[�uA|ĺ�:`��VJ~��0���}V�ʈ�\��Z��|�M�������ux�ϋ�,c^�A.!u�iU+YOW���s&ßy����T��['����T�T(�*���w�aS ENZ�%�TW�c��o�N�h����,6�t赴!xCB�v�?���IIȆ���~\mN��OPDQA�i�Aۏ$-11)��u1(���3{p�1Ķ��V ��'Ԯ���?��dm���Ir":����ZV���
�KW0Ѵ��r���o.�;�1⣷��[yUD��>.)���"6~߭�3Pi���P$�Q���)���o���R��fTWj�g�p8
�>�a}�4�����?-�p�4�WᏮ�+�EtQ@�4d���sT�H-�Z,D������a�­�I�{Й�����\��f�����kx3:��k}���s�A���p���j/�b!�ݎ3��-d�N�iG�e����glcT����W/�Z�5HD�)���^���<$��Sʹ�DK@r�
�,&)1D_��Awk��L���𕙐H��l�<
�@g�E���,��a#�3\��*m�Ih:rgX{�0��<��{pt��`��e�O�a�<�1�v����]U}�v]KRxW恾������31��X��?,�,�k�U	�����˚k�ϒ`;�`�,����hD��Ɗ��BҢ%#-�J)[柲K�BN\P���K}���@����ç4/ԝG�l
��ښ��)���G�U吒7]� ��u�9�Wo]� ��k���oZ�?.^�J{�)}v���]>L͇��h��֠�Vr������H�ZmT2;z_���=Wq�.d9YS�V�	9aR��?]9Df�H���wQ��/Nk���ql0�����B^&��(��4Գ�����')#fe	��(R��f�3�(��rG7�iZ��aؐ�Hd��Ʉx[�}�E��ڌ�iR���]��7ӵL�Ne8�`���(�*���U�����u�-*�������G$u]�x!*�ұ��hж߉�%��w�KҤ�U��h4{8�^˽��J�̚��(�4s����."okT��� F�{�)��t#�
�D'�^{2p��qfA���������nS�'��kR�:�$�e��&/���A��ߍB�QO�͍@�S���a��O#�����l�J�� ��h�hV�;T���������j�[�-����h�y�s'�JA/�Y�!Y��A�U���:?����o���&4W�'�AyY�=0���ٷ{�.G�g[G9�ʠ%�=�_{� �D|^�*�Lz��K�?�P � �<$�w~��7�pU�p�kǅ 2�
�B���F�Q�R�?������Y�-/����F������\���,&w��K� ��ߨ��g�mظ�`Cbe�a9�3����FOC�*G��i���{�l���cR���6I�Xȸ�@Y�!�ЂQ���@�Mr#��Ш��/Q �q@L��R��:H9w��34���J�v��+�������r��?�MB��A�g��v�R��J��|��Խ�4��0i4zO��%��YV��&Hf�O�D98(η �h8	u��U�����؞T�2�}��s�C=��H�֍n�|�#뛄!T���-(��(�l��U�Y����BA���a��K[{:�(OX�C���h��.�ύnN�{R���Mp���H�c���WZ�°-�yI�j'9�l^��P���HݹQ3�C�V9H��]8\�~0�z��K{�cVWo�;���7���#�݀�69���)?V�I$�>,��+�L_��Sr�RC���&�i��^��#_�e?��O��m2I�<_�a1�.Tќ��q]�B��\#�K4U�-���^�u�G��_��Qd!��nbk�WW��&�t8���|�Y==�U�� ��ag.G;_! �@��:�B�Q��<g���&��V]��s��jy0f�O8~gV��a�4�v�`&�p:ْ��8<U�c�;M���*�d����_!)B{zFo���.��J�+�A�q`�d]��u�&�Wn��?��z0v�DR�08�^�I�.��^4�0��1�m(�n�1a�u�F�!LQ������w�_ނ]�k�MXU�*���^�����?�*���6��!μv�@�Y��wE�CA򼸃�pVj�Ք0�+���E;�_��&�"������ITxl�U���8Y�K��%w{X���E�3'G"��Ѣf^��˰��
n��_�]Ռ�[��$�y��$��L��5@Y�\Ѐˬ����/X���0�'���?!M�`�>��x�rkL-��V���Y�3&�Ө Ca-����>�Xi��*B?Iɪp�V`�Wz��$�GR�1�ܩv{�/�[�OY{��@-�s����m�����K�@Ku8��������I-L��f� �h�![��puѽŞ!4�p�ʀ��[�/�l��?*`�d�R�]�Z���#��Q��Ķ�I�
�9��uN�nT"F�Z�ce�U0ʭ�ԛ�a֔ǝ�+]v
�"	Y�&e�h���K�E(�7��U�
��vg�µФ�~�8~.�/�b���)9�8{w�|CÚ&ʦ���e�L�8"��{NQ��BI�z{���.$�I��/J��~P�٥)Jۊi��λ��$.2��j]"�uD8�1j<��fl��u��>���{9<��,|�M�XY�O��FS�̄�m�� v6h��~�VV�-T*�$����cQ�ݭ-�F��w���v���6�]���j,���ơp^�;��=�� ��g�º`WK�wG�%$-�rN}�Dc���8�����r�ĝ�N�\���Ug,