XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:���J���C�8	��j)�ü�2bn=�F�^�T$&�����#�*�u���|��&�aL����i��ÇŞ��G� ,=\ݲ��D;4 #�%w�~8���M�:U3�S4��\��`4J���<<�5%��s��ƩXGޢуjwA\%��S���Ak1��D}D�X\��x`��a=��o�DJ���y�C����L�d�7��w���ќ�)��S���R(+)(@��3Un,�_�(��
�<��r���~���R�T
$q��뵡
�\�;H<�/yJ��@3E��l�V�-�.>g�9��*a��iàĪ���ڍw>G����_l�Ү�0l�Ȕ�1-K!�Y�9��'@:���2XW�0�b�r帛��V;�>Yl�<���Qf��K;7�{�@��U'5_��a��شB��,��<5[�W:��S�{y9�Xi-e+'��N�n�b�KZ�a�]���P.L�ק��\z�l�a�ȩQ�
�V����/O�!�ZE��6c�"}��,�3���!��j�|ǲX��Lnh�|JP5�?"�o�1��H�2�u%��0^'�9;��h!c	`������5�r�kd�&4�wĶ�6m9�*�S�GdF�����$Q��'R��R��X��.�C�WF��F�\��`��E���x���-�����NX�)�(!���]�Nz�&�:�ף������[q��m�%�ӹ0D�y�d4~W31T�ݚ���i��@��WK�뻔 �r���F���XlxVHYEB    500d     be0(�g�J˘�"聂��,]W�Kb��~��;��'�F��J�z*��T�KP��N����CR҇���g��o� ��P�ho�(��.��e9.����ו`L���*��!sw?����g:j�E�����91���#N���|��y�m���P�� \w�Ed*�5hQ���em$Є�m'Tm�Ų�7|+���<S>]��O4�06}B�x�t����+#�a/QE���ٰ�|g�-��4����!��q�c�ݐ����Eb�����i�Ѥ�FEn��;�tO�n�-�Og�$�&YۺB����;��,mz�Y�z9]IH���@�U|5�ck�H�r��Q~mq;���m�q�Ј6���N��C���y����	<Z<Ixa���H��3�3�m���w�jpN4��2�t���:�!���`�䡈�i O�tx�H�,Gx����%�U'����@��������>{f�`�H:'1���E���XK:� 9�DA���H�1�w}eOMQ�v����`�ZYKw��ϵ��~f��-���9D|�"O5���s��W���z�RY#@�>i�R�X���Y�:�����\��أ����V�J��a��k�N� ����N��2�!x5���^9��̱TY�8����<�A�yu?�)c�C�'4Qh�}�[l�>åAE8��ܟ���J���#�r�
����ɈG�k�P���{�Sn�o���:��;Z�hO������knJ��@��,��}��~�x��6ag��;�,1��^fDoF�ܠ`�!���q�:	�_�02�^Y"��8�o��5�w+�����7V<�,�����iS��o-�|s	ŚAي�HqK��[�Z�zbB%6�`:��"z$�h�F%'�$[UB,����(�'n^��dښ���=o�%.;�y�AC�m�}�k8z�^W1��]�������� �Bh���E�,V@<L����/r�9��h���>2�&i�nR����nW��W���{��I�n�I����wI@�\~�>3,����#
%����`}�����<]�P�kw�nu
���~/�#�i��B���¿݊���![����Sq�MJ�68vI`���^-P��ŵ��S�|7����i��:���� ���'}I�8�P���.�'%vd3Ұf6	0�7H����@
�͎�r<>���
:�&Gk�t�a�1������6z-W��s��J����D�V����EV�W�R`5B=MI���0��@�x���J��Xln����"eܑ]���o��
@>J�P^�IDW@X�k0�4�x��P�-뺢6�J�%����U�f@ *�� �dp�?a�����&]@��#��ZV�����PjD>ބ=ƯB	`�#��] 0�nQB�����R�����b�DF�g�{my��9O�B�>������f���h)�����1����;0�P�>���ޅGc�D
�X�-M͞���R�Y$�grd�RZ��@��'�*��� OOv $��H	.!�6!�m��8jܺ�۠��$S,t��k+S�=�����ZbqP���U阠R���^֪
�T��/G�"mW�xIx]<O�,ѥ2ɨ�K9�o������~��]+l��yF4�MR^�S��f�q��ܗK~*p��FX�Q�ba|�4@%3�"�C�����!�w��бG�x#?zJ}e�쓷P<�%��t�%���<�k�b[xV�Jөႜ`;U^�t�cń���F��U�
��XN*�ڜo��\j���	��K��Q�|G�B<����	6�3����u����o �I8s�?R�B�ב;s�S+Jkݞ�������.��j_�F@��)��gH�?'�'�:�A�9�;&���Q��2:�r_Mk���)�����y>����``�Pi����� �������a�2]�F"���o�|a��r��d�
��B��G@Wq@�J��=\�g�n�_��_���8id�#�Sli��Ȍ�RĨo	�Zk��$3�:D���ϣͪm�ì]c�
������|(.A"'tj���с�Q,��id� ����|+�����~����՜�3����D{*^�Yty��خ��:lO�5����{���z|8V9\ol�Ge���_!ߓX�-��S����������Ӌ��7�6e�_���b��U���"��7\{�5 �`(H�5:p�t.���P�	�����N��ް��hX�y���DiG���qu�7���RH\��1�*#����-́��?'��o�{�ّ�(�^�/4G�#Z�f�)�YT�ʜ�����l���c�����D�:�D�0+�ٺ:ZJ�H_r8��x.HN"�8E��K�i��
}��uV�c#Uh���p,,QI�/��xQ�1�ۊ��^0bFꄅh}I
��ً�ZMt��4Fz�����}Kop�Ip�aXV;����,A��_�n�z8I1)I�8Z/�ܟi�����3TQ�p�7A�z\t噌r�n!���T�c�~"O��O�^ �=2���5h�ƅ��!�ZQ�%:sO�L,��k���G�৑�"������V�����[}\��Њ������E��~i���u�&E��?N�y��`��Pw�1|�an������ɤ}a�*�����e�r�"X��APq�}����1;�:���r�;�ږd��t����W�!}�S��93�s�d��[���9��c0�<����8L���h�PN���3���GbFp�-��k�,��-�=l9�~ɇ��b��4(]�@b����b�	V��Uyn��1�]e}��>�3��;���f!��ְ�L4�l���㼭������eip������aV��ׂڏ�X��;����)n��_fI� ��ݰ��0�e�Ȭ2�������齧�rb�� �Ć��y�)�FyH�1��;$9�
woL6`)�,b:�u��o�TIr�� ��