XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g�޽��-k�xԎ�O� '�$��V�-����I�M��v�lSii�7")fF���9��
O;>6�߷K4�2�ǈ���R�r���?�@�¸�h��$}\�H����'�<���e����m{�E�[L��8�)���3�%g^�6*m���A���4�=����2�&��	�ʦC�%cX���M�p��#�o�b���qU_����&E��-����Y����M�l>�� ߝ23��/+�ؑWo
D�-ˑ��<�pxr5�v���d��q�Q��Bh��y�=L^���?C�q��P�7a�4?ܱv��҄���$%I�tBA��S�>@(E�����{-�Oi�-��o�J������2���Y=f=�*�ցJ:�}HG�g��ž:ɁW�%�XIHҢ,�j������W�̭��I��g�`�hgrt�O�Qɻ���K��o�I�f+��i=�n[�ڒ{*Ƭ.���n9#ll���#���`��y!p=?Y ��/��]��$I�Q9c~^�lIas��J�s���5C�@��t�������$��(�n�U�G�X-���h����#���֟�r�h���0婥_�P��JC3ll���[.�G�Wt��Xw�E�n�u2֟�ۭ>#"_Yd�T*f�7�k����(]pkH�^�J���ۥ���yB�O}%n����^ �6g����ӋByf�:�H�b�d5���,�W�;}v��4iCHay�ٌ��c�����AU�'d��XlxVHYEB     634     2506��L�����h���2ɬ �f�&27��E�j�.6B�/��5$T�P����׽]���06�]P=caF
��m��ޔ�E�{&����2�}3�hp���4��W ��?:&;�[�j)�� ���6U���N��}��c��-���ʷ,�/�rY*H)�ů�����S�TpRW�ׄgp����H����7���M�����5��@����E��C%i_�hU��o�${��$�ALK�@[>D$y���A���?k>ÂH0I����k��\bͣ����K����@n�k��ܭNKY�8�~�$��Ou���[�-���E��z����g�V���_іA����4C;f=��ɥ6w9�C:�d��/��c����k�gNgis�G��v�鏲�^��v��~1��)�$bd�f��G��H�/�. ����M��Dw /��#>��/ PR�H�ϡ���N�bD2"����R��=��klT^N�J_���R���$�_%]&��p�6��:,�	�w~����ֶc���M뻤h���u=��V㯑k���$���5Q��������+A�$n���{dcr���[�