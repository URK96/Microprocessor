XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Nd:6�� ��D�����������KP��e�&�Έ�����>3�����@���<�)׫v}X=���l��EtN 4�/�W*S[]կ�v���]�̲��m�[����d<j�����=A�����B���m;�t��n��!������s%�4h���-o��պb�=w�G��S<�$�J�EG"ڥ>\D}��f�^�cDL~*�
�PgY�ъh}�s8���cHA�A61�o���ۙ36+�X��eLBkZ�H�GL/��E���f�N�_۹�bj(NYU`�G�"��r���f�n��r84�{;t���.�c�?�$�]M�"�Y�\�K����wJl���M��w�NM�K�'>�K�F�S��p���N��wE����S���vp�e��2�u"��,̅�Ly�t�4|�W��M��g�e�ޅ+�g*s��U4���� g@���Wx�:p�Z���IEFlCB����P��R_�ˑ�Xr���{�vU��	U���B��}v`��ck10�`���~��͔����hm2�� �,'�_��F~�h�y�?�05���_�;JT�[���b�r?}�{	 b��15��^F5 
.���ui��i�҄f�����L�C�:��/�70+�T5�R�� �j�K�v�{-\Ŋ�\m�~N�}0gW���Y�_��bI�ג�>����仰-G�$�9�|J�C�KU���&�u�|c*}c�ڽ6?ɱ���k�Jw�T��ߣ:Q�H�c�����ͣ1�W|y�zXlxVHYEB    10ff     490
$����V6������]�p��ؓڇ#$��>�� N��aѰ�q��g�Ż>�Uͅ���Q�8Vtڵ&䆒�MZ�}*�Mo,j.��t��	E����P�X_"����'�	����,�����mh����N���/�Md�p�G���*��v� [�$A��\�͛%��#��Vz�|�޲�é���G�7l@5�j@�� V��P�
!ݲ�������ˬ�g�22�W�`��1�'Fb���n`�h[ʉ�=�淋�����.��s@��'5P�~Y��zM�|���گ���s$nW�@�0��\�e0|�9G�3�V�k�����2��m6��~��h����ݩ'����A�����f��[��8&,UG�6I�/8&�x�Lu]�;s1�������<"'������?h�>M�a���:�E��Ċ�:��:��Xk�\�;~��z�L��,t�@s^�!^p>v=�9V��qxwƔ�vDc0��|��Ϗ�%iֱ�{A��tw���~����$#��9�[r��,ݗ��Q�W*�W��be����#�:�`�1��.7�J��)�BS�ܒ4��;I"la8�9đ�;ƿ7���gq�g����%$`��B��^��1߄�����_&���Z��~��'������~���p����X4#3v#]{��׵�G��l�t ����AD�Zߘ�!���Qi�n9q�������1��01+<(m����N�����
���1s�����E����bױ�j�oS�]*A/H;%�
�`䖥�Da�#�.}���8�����6�wTO���E����f1�����?8C4�oA��o�������w#/ Yf��Z�l�
�Nl�}�+�]D�� �fs�u��x�����IN�y���na�@������IB3�ǳ�Ņ2 ��3�F:|��|�G8�!�m'5b!f�DV�9�xOBv�tՖ��!x�(ؐn�*a0��p\0�$��'��g�ٍ�/㹺6����s�5�y�P%�v���q�-������/��8UJyY�.a��hl/Br�;��G�iQ�|96Vr+@|�|I%�8CYP�_�T�wʆ���-V0>b�t7J�uU4@Epr��E����P���ʴ�gl��ΠQ�N�xa_jM����w �b