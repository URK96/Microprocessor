XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��U*�ݺC�L$��S�Bo�XU��/z����Wp�I<�����P�k+c�-��_����r��7X���j��2�Gp���f��?H�9�o]�#�Ğ������|W���I��j;�u@��zDkCK3X�������~x��l��=w*%G}�8޲W0��Y�:]���ـ0�p8@w�w&�� @]�,��4c!|��P���[(� >�EG����	�i��O!�WS_|�4�k�"�17�6�i�c��~+^�����4)��ʊ�����km"���8ԣ��G%)���+��3�Bٯ������Z��P��a?����H��9���ނ�Wʾe~VH'�k�6�}��k3������ �Z#�lȰ3Kf��2��-XT��B�N�el^5�3	۝��?I�Խs�E���Q��jo��HY6v����/�f�d��ĔJ�m� L�_�:��:��O c?]p9}��I/��X�'�����R�H��G>����J�|d��sT��[!.�\�������X\���8��cA��a���w��*x��%���я��N>��Fb+���+?̱Xb�7���58ס���X�rrYp���ڦ������� \���!J�~;LU �>��\��w�J�#�����p��3�VMk�=�TU
�;F��{�PL��n �9f�������t���7�E2ȳZk�Nc���ݬc_#�8%�p�/���Pd�^���1J��_��'�a~5��:�+�xXlxVHYEB    41b6     c40�L�|Ux�H�Y'��z�g_�^�D�U`=nFԂ_I����imo/���A��LX⪱�E	�:qn��sa�R �Հ�Xʬz0/l�ܷu��v�۞��7b���>�:����~�]�D�E��HsZUTɞ㍙�E֥(2�a!��|z=Ts� �g ���;^J�h��Q�s���T���5� gO筻�U�
2�w�}��]OQ����)�m��2i���>��nc;��� �lm$��)l�BM�I��7��I7��9=r��V��G���L����H<�/�͛�q�[XիT�CG����0�Vr�ᲦAg���g;E�ʁ��ֶ�B���Lu}j��}@\�d�Ʀ�r=]��
�lM����y��E/0YX�J �s�7�W��"��nn�ݥY_��i���b��YC������f����a���ɷ�R�^�ݞ�L����f{Ê��Lz0gw�~��Wk�.V$ϰ�n�ܣ!�#R�Ҥ��QA�㓼�xQ��C���]%��ɪ�*�K�,����f��Z��v`�� �<�3��2��"�O��|k��6�����!<R�i�6�U�5��f�e���\��4�I����L9�A@�{r�n�����4����m&:)�	����*�Z5]>���'��M�����s1�q��כ]ML���`h�y��W�j���'��c�����~�d�A$�<V=������:d�h1(�h��M=*\�\�@"��)����h$��ݔ]��*��^��`!�x+,�����O��X�%H. �����\X�u���̲1�.2�'e�b��(���N��G&�cr�24jj�sR��w<Ԑ|!�M99˂+���
���n�
�L�R��rd6a��>�O=�,��;Ւ�)
�=�:t�p��Y�tI&�.�<��{�@���h	*��}�.�W�kr�F�G=��8P�qsi�%�h����%�Q�g��z�<�3����� ;G��?Le6X�k�S���a�MsR������&����7r�����H��u���+%u�v��A�t��fi\u�R;o7�?"B�HX�xH 0<�i�4+S�3���)�����	�}��4͎geY#����*0��k�}t�!�齤h3�X�f� }O�`քv�)^�Y7?(��qf��	;{?���[~3+ΔF�5��#����q"335ٶ<0�;�F�\�W��k�:]|(Ӛl���\�~�7O�݀�i��3(���!U۠#J��avp�B�	՚��I�o!3qu������c^�(���<����rP��M�P��VeI��t�C	�"=\��AB�Y�``7I'�kO�e� ^Ĥ��K��z��} A�.6�%P�S�$w�[��bÌ1[-� �@��1��M��́|��u^�Oz�>'��j펬)��C&d�]�5�N�Z�/4�gKz4B:%�m�D-�Ω�z�#&��*�1������ �~�� �[*��|��	���_��O�gu������rQl�ԧ>v'T���9,_ȳ50��9�2���էk�ԉ^5�nQO͹o���^B��_\I i��g�.܆6��|bK�P�譃@��w��_��F7��U��]I�����<Le��ˇ����)�ߧE
kH��e�4�nX�z�TjP� U������)ش���=�}���Șt4�~
�0Ŋ�#�����>�\�h���EN��0E��Mg�B2����3�2Bf��Qdo��(��#b�m�O���0-��om��RI�1i�n��a;���G>��ܷ��oLg+�mKe�6�;+a�Tz@��uIq��WT��\�5֎W��y�D��!��y��9W�#ɫ���&��,����6VM�R��E�x��v�n�UČ���W�.�!���켹��X�GVE���<������D��	b$�y��$��wr�B���8p��B!�ŉ��a+&�'��7i𮊚0v�e���-����;6�P�����]�����zwL�%V��K*d�>sC�C��+���<s9|����&��e�K�J�j���f9 ��cJ�'�����N���a�NxIRpd�s9�Ũ�T��RO�p�}��ٳH&?@��O2Ӏ�6ۊXPR ��8�F�Y���\�J�v믂U�@�9"��K���y_2Φ����������0��A�Iiw�,�FX�\	���)g�sM�ł�7����]kF���f�j�0�:��Ͻ���
��jɋV�����ɮV�߭�jP"���$<3놽�=_φ��.��P��3��������������ʪB�(��?tgE�O��L��%��94��f��짷
�Za_��F�P�
���f雪�p��w��ڳB�9��"�ZC8^λv ��;�<�y���^ �.L�r�g)6"�}G��{��Y��C	�&�5dq%o.G� ��m�",��?FFN�m�!��d��F�)�%=���r��fI�~ܾ�Ƣ�"ߗ.���d
�E�c"+K�DH ����̀6-�{c@��ޠ��C�[��Ʋ�k���M�߀��q��T㧋�J�R~z#U�)��r���U�Ƣ�P(z؏Æs�}���U���a�齋P�v�o3����go$[�s0���ql���y5$��Kv�^��XL9�V�1���l�/|���\�N2��V|��'� 	ԉ��/��r��7��YU�@I>N����4Ȫ
��->�#�9!L�z�BV>]�]hs�M���ͧJW�LWD{�/jgw�����d�[�7��m[xfg
�u{�A�\n�Q�Y�۾���å��@��j]�0t�E����)���h^��tQ�b��� 
�&?�p>ϻŪmO\:r�Z�N�N+K����aO?[�`�9������m��e�T�`����:�b�&WawAs�/L���/=��r��9��'$ �dK �˼��H&u�u�<��"�r���^$�/4���~��T��d�J��&��Zv���x��jN=�AD�0��l�ϯ���:�b�� S3/ޢ;����\�r�w)[-�އ�aoBV�r���C�*c�g�u[l