XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��L�*�l/d�	��\X���Xf��V
��ؘ<B逤�Ѕ[	u��1�M����x����sw�괭C�kz��3|�	�Ɨ�\V$1�����g�'�n��z[��ܼ�^���6�j$��##�9� R�`��������"��8�dJ�d�j��5RyKػ�1-���q`��s��m��s�N����fA�����TPG]�ߨ��Uy/��|��Ҵ���H�v� �mv(3�u�M#I�M�2Jϫ=��$�)�(VXȯ���2��DK���^]!U�$oj�~��h3ot ��!Y�4����=�
i����"��!��s&�&6Ԏl���띡k��ks��>��Y�o������F����
��^���5D����@cy���f{�a��	������Ȳ\��x����e�A���Qh7^�H��e�
;mǈ
P_�q_L>U�'����}H����Ռ���u;_�%�$$����{(�6����j��s��H 1{'�U�˄�t�U/@&}��r�P�Mo���F��B��~SD�SӺWN�xȗ�ݺ��
	Q��='��zP`4{�#0.*�h>����^\�i��=N/2�BQJ%M��6g�V�B:�L�������]"�@-`-4��,6ls��Y\��>���{� ��"B�9~�M�k�u&8�
�;u�t塞� 6����K�9�����d\�Mȴ���9`�#*$�
�i]E���}��XlxVHYEB    41cf     c40��K�y�a�>�z^L|���,�	��PG��n��h�Y�bU$��O�*4�Op8����m�H�{\B4I2��L�[��0�����R����@�{�4Wv�O�q�>���㮶ՙ.��6�5���	X��C����D�Gר�.��sH���Φ�\��d5|�^�_�����Դܢ?��Q'�-&�J�j-䕐�[��>�bQ<p7l;�����E�>G�a~�lj-)�����HBQ5��h,�l�2%$�}s������ZC�b���'�̳z(��^�|�E�G#o�\��&):w�Cp1L�.KE�M���Π��hs�	��-~K���Wd,uI&�IϘ}d�.Q��ۿ��.g��;QNg��ο���{[�9n/��Ԇ��p���9�EYR4��)���3�-���H���+Z*�_���,�o�@�
Ao��oԸ��I0�!�d�.Vh��Hzh*�;��k��zxԣeeic	��#���&�.��?٭E���ݺ�v� �:q4�~�z�ߧw\�/H?M�ْå�m?�,��u���\��CK�9�|E����]�Ďo(��zy:�������nC��ӯ�?�+##����j7� �q*�&�r����s�|��.+�旯�OV�(���_��Y���|�|!�`Y^84��H����E�,Ԟ��g.�=
�߶�u�9)p�3�+6�0�>�L|}�e!ZV*��O���a>�������1)`J�g��d��ޓA6�B��� 3�-��$:=߅B����5���EkSC�}��i`�\y���#~/����E3-���J)�7/e��� ���75C�ԃ�[}��U�N͊f#��������`�--b�K`�λVJ�����T�,Bc�H���d�`�T![�@0x���.ĵP}��}��Q��*�3��-� �ո*]px���Jȭ�ltx�"*}��ɵV�m��V���UҼ�#����Y�HI�_�e1�O4t �lN��]���Q����7rC�|���2��cqU1GdU�qn���6��R\�Ɩtz��<���╀+�l�x���������~ȷn��İ\>|��)�.db��m3��a@��%�ᚌqoL��p5�=�nk�ZOm�Ch��W��hh^�tc���F��\����%�g���N���\Ө_]Uv$c�63u�
Vl�<R��s.B���V�!uZ5��Ñ9Q�\C�+D���=�`�l/�=�&�O fԽ��F�W"4'b�ʗ>鼛�B���>���Ӌ�'P����]�H�,�ׂһK#��}�`F�c���E�?ˎ��P8V����Q6b����2FU�{��&��@5m�K�K�zw�	4m��".
�F��p�*��
�<�5)F�$��g9}�~"S��P�&�q��j�D��GA�:�(ؿn7fzo��c�nn]�|�c���\<)�!�����s�y�Q����}m�gk�U���~���>���A�@�[�J0�~�i$u�o�S�v������T|�Ơ��\]�R�ʭ.wh������)���6m�-�>KKd�����C��T��
>�3�،���e+�e����MH3Q�Hk���H���O\(��Gƹn}ޟ��x*�C�����'+&կ-�.��Q�x��>z��'���+�
�t���E���G��996�g�CȦ��?��9>�;��w����A6~Cm8�¹�� V^��~�����]�5�_�םq{M���h��Ïŀm�q(@D��0�# ��SW7o�t� ��Pl,���j�j���voZثH�pQR鮶��m�αd0���7(p�D�^P���9l6d~7�������ui�ć���9��4At�&�$�P�������zz XS�Ke!����,��D@��M:�S�\ք!�Љ1y�I���g����#��xS�Ȏ�-c�oZ�l�E9�D�/�.:�a��eY�;�~=�W��0ߕ�UD��@G�5o�i,� ��`
ƿ	����iF�*6�D疰�e2I;��fX;�t��m��n)xb|�g�����ղoԿQ�iK�2�E���xa&���Q��A|�I:ͧ�4(�c��VbG͜-�W�+� �$�`Cu�o����9�:�Gfbdݡ�h �5}W�zo�KH^a��]�3V�Vs^?�c�ʽ+pk�9N�1��<�	������+�eW(P>�$��I)�1�ɲ��<�V'�헀��?�5c&e�d�y��5��a�O�30�	^VG�0r���ۄ����0�6Q3���ʛ�ւm�7�%9��@*������ؽa��_s�[bcQ@[���K[̤_�m"��=y��'+�͕���ށ���=YxE鈂��3\r�Sd�
�ߪ���1 :�i�U9M���H��0w�<|��_��y;&F��&6�;�ǧ2���?&��+丏8v��
 ��K4��A�y�W�`r���,?�I\�p�yNFSE%��~��,���Q�	�>�Z�t���N�Oȭ��C��(8_T�}��,�n[�NL~�՜/Htu��ɎV��T�4��:���՟����.��^f����qǎ#�Qg�5E���-�$�d'��I����5���6q�֎������0H�����-S�B�@c"b��H�P�񯃔���hd����̉` )D�A�2�D���s"��T{�b<��D�Dx-��Z,��I�'~y����BH�Ŀ�6Y�b}-F+���p�ǎ�����*$2���*���Y��#1EnJ�{!y��!F����bm �$6��A�^_HΆ�@1G���;XK��fΪV�������&��XD��������Z�:�IB
{]��ܑ%�h�;%R���9�Z��Qs���&�
k�Y���I�Q�y�\25�u�b<��L��d
{��C��	h/T;���l5�,�
��]� �����\[�c�^�'�ӂ�!ZK{>�qA�����ޚ�7d� a��^�Jjpa^"�,����0�d�^���,%���d���or�����/���w�D����iA�j����� :p���Ǘ�u�.>n,b����I����$��