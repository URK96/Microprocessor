XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����E纓VAi��qf�����UhG4L��Y���Qp�����i��8j���]+�h���}ʣ���[��9&��?��\�\Ȉ*�IG�;��.�2��N7��|����]�-����)W3�Mn7���M�����ɧI�̍f1�QF>���eC{<Z~y�4��f�u�z�a�Ì��n~���~r��85�4���3&3��	8�6hD��ޅ���E.����=�ry�璓D#�81A��m�EB���(ƒ�$q�:�e��D!rao3L�j���Z{��P��i���N���W<u�Es�}�O���?� ���p���$ϣ��֍����4T��%vm�`���a��b��j��5>74���X���E��z�+�0:�e���!k+H�:��q}�h2M�kb�I���5 9��/��X�v��~~OU=�.P:Mx�غ��`;?�_k������m(3���J�k~r��9d���7}Z��E\/
Ū�&�o�y���"�T.��c�ǬltD�DY@ Í7^�i�B�D��%��8*��2��'�j���t7�AB
����V/0��<��,��&y�1�ǌ|^L���WC�aF��;<;ڌ�5+����������Y񿮁(����}9�ވ�@A���=[��oXD��>/,�Di��ؾŜ$'H��J����B�l��ټ�4�9B2У�+�n&�Ok�����O{�Xܫ%>�.䍤���u��3S�)��.:������`�����BXlxVHYEB    edab    1ad0)�אuL+�s6�d�c�	k~���Np�^�3�_�����.忶�����9�[�Uo��\۳��������o�����Qߐ��u�d0g�m\�m��Π����4�-�;�J�7O�y#�N7�*L�%�N1T;�0�f,X����y�0 5��2:ZJ6�S.�cg/Ce��	������X�os���Δb:�o�;�\7̾x:�Dn��sp��ְm�9j$�dCZ���ꅡ\�3�~T����.���1@�nC��_V�Z��% �U�M�rLY�G�N?t&���GEMy{-c�鬻��1�v�x� �>���dT�X>����R#��޸5���cq� �#�[ѷn+���׶��){������Q��@hz���	P�,�M�j���C����`�:���6�C����F!78$�W���;=OAÖ��NΛ��q��u(և<��v�X�pQ<�bw<EjP*���ý��o^"��5�n,��J`1��ۛR��\���m]�թ,����7��*PO]C��}��@���/[��8��`܎o��!��!z���N"�����R1�H)su7��hJyK>lJ�ᗳu���3�K7��/�Z �Y0�����Mj�a�=tvH��L�%�����V��:@~�#����&s�����)�� 5��fU�\>r}�s�m�OixL��#G�̖��GQO���^q��Sw���?�p?�0�u��t!���� D.�琄����g������k�(N>�H�Nn�rt��ߔ��r��ۙ�Q���Y�χ|�tQJZ���X꭭ZS'�\�@.'!i����e�mɵ�r:Ժ�;S�5ݥ$����"+���<���?�Y�T�V	�8�60�C�BR��"�����7E�
��z�}��,$T��0\`�YF�H�ʫ;:.���@Q�"+ ������ y���O�X�uW$����m/w<�ܱ>�Ĕ�0�.,)C)��=��T�_G<z��0��.B4���P����#օ\e�
���{��y�����z"��������¡��-]�:��tL�)��cZ�'&.�{�R8m�����5��K>�����p��!,ܥi*��� �G��n�y�l߁�ƴ�.ӊ�����
��?��e�n'�Tzku���۠ۂ.���	�㽾��_,Ca��-��9�7}Q|u{^~���Y���,@��V����<�k�[к�'k�<�s��|�|q�@Ѷ��-�s��_��
�'�����tҒf��)i|�@�f!gЏPD4�-I@p'��q}1�=ٳY��8I ʇ��4OS���;��y�����	uܪ5��!�&E闋&U��G�u�o�F���S��R�K�cu|�+mr� �| �,�e^�	l�Bc��(����Co0�z������9��[�}�����.���{�]cr�/�v]J2��T��>h�~HܬN�����{����tj6~wq�g�fp �Sޯ�8��^0�{������Ғ3%k�s�	��h�{l)<�K9�	s^m��4��f{�U�����,eJjb��#��}T����T�i��@�["[�:6dKn�*2��Z�Ķ�����Q�'87��������j��Ͼ���}Br����C��x4f���D�׳�5�QR,I?G�� x˵�El�����r�`�/{]�3F�+Ө�ly�$ͻ�ը�r���}�^Ѩ����@>[�U���>%(����_a�==/(���M��3�p�q�H�2��VQ����f���?+��F"틩4��J��,ǐq��R�˹���im8�\�+��r���=7Ŗe��)��tsQ}�P���K��ɴÄœ��S�����c�:�-���^I�8�6��V7�lI��x���{���^F\ƽ,@�9�h�>�)�]���	)<F�x�o�C\�-�9q	KMD�]0�u�MyR`��_��Cw�8���p�{aqҪ^���z�PC8�1�Fb��~��h�no�$[[������mVcK�O:��S-���͉q��o�)�,���N��Z��rN�ňi|ks1�3���Y!(F����!�����n�r-�͞$�l�N&��I�ᛀ�I
���kQ6��A>ḛ�Bߡ�%�G�c��A �󷁧*��3��l�K�9ы�lj��oN�Q�l��p[!�n��L-2>`��]��_;���]����,��@];R����fR߃_�l�� � !R�C������܉����"�����yU0�+�pEnħ�~S�A�(;��E�#U���Ƴj���{߳X=ꂳ�v�5w�Yd&ma���GE��dMB_d��5D��*��<¡�l(P9o��P����ޯ`��ҼW�����t����.���[P�zrO�J��N����[�`�=��Q|ée��E�H�臐�_����=�q���_*F��j?1B{t�Y�uE��ʞNT��2D�����P�#��S�hB��f5�I��T�V�+���I~א�P�hYп���"!*�\ Ǿ�ۘ%O�.���Lf�G��u�����C;]P��b-�>�G�		�����k��N����զAzG�vS� �����6�ÊȂ1��z��eН6��k�9�8�8�՚�p欍0�*
@>���y������O|�X���ص�a�-� ��5jD��O�%�v5�r��l�8�����g
�7�޷8��a��x����v���u$E��w,�	���+�!آ��=7�>[�ϒ�]:U�H���5�ğ�7�������8��3݋���W�v��Ƙ��;^q ��"5��"�Ҟ!Er~���RV-�2l��Y@Kc-��!��m�\�Sbz<�.��>�T���
H%�S.�^6b��[���p"���k٠ճC�5;����2���K �O��@�O#���޺��!�$����)��R���)#�m�"R6����o��r�pgH��GG�U4��,�눧�d5֭I�_�1��oc����p��ָ�ꅓ�U|@!�� %f�S��tܰB|��C(�[H~�?z��ߛ�$^t0]S�6��W��t9\?�'R牕`ߩ3&�;��6j���4n,)�`+	�6�{���K���4dGq�>,Nɴ�f�\="��;�H"9�N��N��Tߢ�������A�G/&I(�i�������̸��v�4I���&]�
a��W�d�r�KP�e*H3(E^<��������|S���]%i`�������k��k��}C�i�.Տ���ć��#��q�N�=v/
e,~c�1PM��7�'g~4o�=i�<i��ħ1���k5P85!�����>�]�@��z��͑P��,0��5�{`�H)���4T�!�OR�S�N��P����l�{�\E-a��������ݵ3j����"j���E�k��w�zꑃ��4-�^�)�>����,K�u��*�eq�.�Ж�S"���UB������i
�OE�0�� U�PGn�V pGr5?ԏ\}ܓ}HK���"M$�i��Фg͞=�3M{1d`���ƇL�qf��@zYk��#��'Kԁ7!h�|�n-R�����'I��[v�N�2v�Fn����!9#$픟���tDӻ[G�9E�Y*:0$��@E&\�*�h��qC�曁����PM>(
O�M;��U��5�6�Kj,�,�H-��E~�*ځ<�ʺ}����|�dYF1��P�8���O��wK��<<9�ҕ����g2����t z�+ǿ#�wS�f��?g~�{��w]%�s�+rН�ͫOm?�k~oÐ�N�@��aD����w���PޅW���v,>� `m��)�$2���7�9���/M���-I���b5�f��x�ͼ42���N���ҙ)}#�"]-��vA ��/��T�oUL3�!32ڂ<p�}s�-ωUfQ�x�Zo%r��t���7��s�����V&��Q��	_��Q������<���K�W"��px"?�c\��oH����)T���A�w��F����,n4����;�.���;Y>`:)����G�̯�5�/��^tME����Y ��"�m��N4��ɭ��p�	�����,����[Dφ��@��5�:d/�G(R�|!l3M�a�R�c+�Xζ���."`o�^"t�0��2�D�Ѩ`�I�R��;D�����0[�i�M�
����9�f���^�ۄ������� ���%��r��v_-��n�N{�!D�x�Th)���>��*G�Ln�:"+��g:�f�W��b��D�7m_T

�{�3���&�H��DB�+Q����	���h񶉓�.{��?�
'gF���]K�J����lO�DS��hx4)�Q,1tV;�`�k���¼Zh��)����ۈ��.>L�	�����ZrK���N������K��Z��-��gM��o��+��/hTT��J��
Ə��>K���
��R���:��-�|��A����}�ä>/���h��#��#w�g�(x�:2��Pn�ؤ��b�ٜ�O���]�/�.�՗X':��@�RZ%m�yC��kJD&�%�*$S}|ŝ��.N�m�o��v��V�Zƚv�O_!�_��Ͻ�I2�ym
y��{�D<�v�K�B����2�-��Z`�}�L��Z�Qc7H������4F�k',w��9��n�X�@�A[/�`{5K�/,���%Ħ����p������[lD�^��ߘ ��гc⒇�u+���S�1f��l�@bm��p�)D��������C�巉�t�FyJk���G�:���'��_v1�ge�ťG�1P���?8�/��~jaZW(}| c�"`��V�+i?ݏJ*�K���v�1�{e��HRmq�T����3�N�-*��3�d�M<�Q �E�Nvv�\�jxKaχ�*���R��X��h�+F�eR��HQ�%/C�~�3܈?kȺ߉)�������>�������hH≙ �]�̧�<��Q��l!'�����.�֠�uGY"I�I��c��ߙ��u4I���E{�%�����E7]%ήb�k��$u,�����:��d�q�O�r�Z�16�[C�����_���O���PB���׬�'��xQ����e��]0;��"{6�|g��(��p�V�ȵ�k��$NHEOUt/7�!�-�5:9���Sp�S���j�stc$9�,���'(���j8s�'�֥�e�r��Ɠɨ=F�E]5���Vφ�m���}������I�,��Kҝ��X߬��jF�J��	�ʀ�r�d�`���;�~c����Y
�R�f�"PKx�Z0s�b�	��}�ZD/���BW��Ǩ���:�䩋Vu�K�M҆�݂8�����gx��d�e�Q�^"��9lF.�t��J�~���!qJG��k�3�����ef�C�_k����t	2�km�<_��"�f
�ph��ё��ź;
�`t]H���ot޾�fB�����B:xޯ�o�����U|��()#��$�E�O,�0j���]ԾL�Ư��6�Y3�L�$����R���@א?�C|��9~����K#=f���;��p_��z�C�{;L�y�&�;�� [���vkr��6����:}�~a��z<W��?�*��l5ٶ͗��N�;��R�7�l��w��Wǡ��X�'{I$���;=9��������-Ќ� %����.�{��!�ε�_TMV!,q��I�,����i�	�I����2V����/.����Y"�K&��aO�����]OZ��-���1ɤvü����{�U�W��y�!oLyA+�a�g��X�c�~@��)���S��4]AN���-Ψ*�ν�|�]5�[Bo�_>�V��)�՞3��w���pR��1_K�}�j�!oX 9��~c�:<�5sϥVO�4��ݨT�6�z���\�\^��7���"%�Џ��-�j��M��L�tiA��8���.�;�O�:>MM����IN�^������=�鲈1`�I`�63{<�4���q���>g�F�P��NMV��X1򾍴$G��U��@>}�=*"�M����Ⱥ�L_"Ԥ汈�m����^+g���L���������8lZ�N���d,����0(Q+�����||���l(;h;�)+R˝�2(�cP��3��T�"ue����bG�|��>�c+�Py*�:���D�� ���Byz)샗>�gR�˶F�����"ku�C.t���چK`m)�$GTX�����,,FcE�騌�_���?x��i��陮�N�G�Np��5�- �L���EKf��	�H[K��cj����f��;cl�\�i��vo�ܼf߾�ʆ?����BGe�9��|M�����DlI�ԭhg�B���ב��8]'��x��WՀͺ�O?,3G�^Ǣ��m�R���y�9�ӃHV�3M�w�y}KZp���1�4@O\�z�'u�WM\��ST�h��H�ga�')��
zՍ�����o/��,O���%��Ms6A��{�c�I�	v�`� x�j���$�rN�{�Y�o�ݖӴ)��#�Xcu� ���q���<��ܺv�⾂�F���0��+�2����.��Ď?X� w��cx��S�S��C 0�n��,>�j�9��A�1�y�>X1.r�h/�.�Z\'�� �}iØܔ���Eھfŏmmº �c��c���tnS���#k����*����PȠ����8y�=f��.�gQU����P�