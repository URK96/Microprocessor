XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����I=r;�n�z�C%
�����6ވ��5Um��i�l��*����	fǒt�e���/��j�N��R�@�U AE
�+B��LXF ����h�3 ��Fc�i�N�e�B.1��`& f/z���=u;�K��w<H?%���!D��,�g�j"�p��p۝:�wn�޽Y���f�5F�R��	!]��.�;�Fi|K���)�Qc( 4������#oKY���1��<���w�K��X����R[�K��B�^�S�g+�[~ڀ�?�wa\q���FOg�nJ褡k�\;�X�A.?�nb�'�4Xǅ�m#yYS`7R�S|�T�5��&��%���:P�y�ᗍ��Z��q7m�q�������d���}Cx �ъ��"b� � �@�MR�`����J %��
��`����'i�M��`*?J8�C�]�hcV�B��;-���U�/��7U'�B���C[G����0v6��͝�(����+�?��^�M7�n�)J���j��?RwY��d�{c���ۀs�%�k���KC�K�j���Z0��G��ܪ��;w؈�i.*�R���ԫ�趨l�$Xz��@��;����C��:�mu��/����ϭ�3��G�J-�?��SA_�w�����L�X
gm� o�񄉇�2X�0,A��f�>�Y\�}~�V���c��Ѓ�^I�J��U�Zn�H�$i�3��\~(�=mG��NY�TS���tS��;LN�yU���#.MSD_�[�XlxVHYEB     6c5     300�&���.�{ ]��W���:�)�9��� ��� �$�8�:�
 >�@���"Q�G��j���H�}Fr�oQ�S�<��{�,�'ʏq=��X���l����[G^�k��5����е��x^�!`(�o���h:Q+R�.��٘41��.� E�7�-	h�DM�� �â�1S������N_@������ļ]vvM]^_�N3�_���o�#�[ɦ��<��?���>��K�o�e����>�����d���k3��>��(v2�G7'�f�L���G�����c+�Q��ҙ��!��'�"�;�	ݔ*q�W�Z;|F���f���eR����썸� ���5��R��eA���<u2�"�h�q�4�i]�c�S]��,� ���T`�K+���k�!]d%��ob$z����'?�h3�c;�Ɩ��B��O1NV��﫭��?�6�離�oN���Ҝ�?�b�6RL�}�6^� �?�=�_{�4S�����-��l�S�O�h{�`�U�ǟ5̒�_R�����^A�(Z?�M����0l�ɭ6�o�;��=��|q_S����O�4�
� 
!^�V#���� , _G��z<i�	3l���E2���Rɪ��W��{i��nǷ�[��y9�(h��
�yEB)N%T�]ǚ�������)U�cHh��3��#�;��r^����(�*qR�q����y��l����4NU�#�J�G ��7�͘{��;���(�n�*��`7%�2�a��y�