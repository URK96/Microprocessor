XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&0��$��{�Q�L� ���W��5lw�!qL.����} ��C����"�q���~ܷ�	D��8FB��������ܾY5��OΦ�4�ͺ�sS:@Z&�/�p��B�t;��y��C��~�جw��=Ƀ[�!Z�*뎲�d�uU�=^*E�lv��!��F�������;'�@8���%�L�}i���R�8חVћ*#��m����헴���R1#��^�K���"kq�	:h�M���,�xz� �S:3�������U�U�q7�ˉ�-mRw˳��-��Д#�1��p��;�{b6���"��O��"�9�����=U��/�w�Fr����4�0�a����aZ����V�H<�};��*�Y���<����2\�B�L�1��t��(s��c���]V�s���KZ��
rً\���~�1 �n�yM.޻�Nl�9�K<i��"� R�Ɨ�@�$p�cm������9�:Q��T��/��Ëu�*_�����2���~�z{cU�)+��AWRcF_�(�)��BĤ��]�W����k�LǆS�O�R,�յ�n������z6�5�B�x�ȬJ���a#;�D��9��
9�q�g4E�pS3�����������;5ݚ�{�Af��T�uB���%Ĉ�3,�{~ʉ$��=��+���8�`��ڈ����(5�D�]���H}�(Fl�b9C=q��D���вܑ�D'���Ua�� ��������I;���D�Ԛ�ˬ��/Ϸ�x��7oXlxVHYEB    9b67     f50	���q�Jg������ӛu��hZk�����3����¶y��윊���X�C��=1���"�[�sV�|8�q���TF�����k"�<��8)�;+}�C{
�Zs�~��&����Ȯ���)?kl�~#PW	&T�4Z��DzF��%�Qt�%�聜{���JLd�e��C��'z� �����+��2�����t,?|(q��{s�ߴ�����
�?镢����P�	О0 {m7���}q&G���1Wh<�=�I�p��·!^������s��������c��_�Ҽam�^�r��D�py�ko�<����
��%�tK�H�͚@��Mt�^*iZ�Z�V�m���KN�n��́�"�Y&� yd��[�;M�O��t� @��:S���|4u�3��s>`�0��u�O>'3���ے;��<�����ɽtqq�5u@����ܭ�"[!D����#E*���i��94]�-]�	������Ձ��^?��l&�f��B���Cx�� @�]�|;9�TUp�-+(�h�BW]hb�{.є�ׄ�f�n�W���
�r�V���U`v���4�:ݼ�B&�vp����fk2�4���9�7E#*�R���)xFz�,�2K����f=��_ u������c�]X����\J��;��Pw��#"VL 
+A�*@]V+�q��h�u��~8v����ԯ���O��m��WC�D�)F�/�P�Ai+`7�9k������VU�ĶA���}
��?ӕT�q�;�]<��Kˢ��8$T�yt �!c���F��������C=��9Ȕ3D�c�v���̄�CmYe�{�y��x��q�x ��Px|.��0��`x�;�Z��[����q�\#�P�������� �)�WUS��lyZ� ƅn(�U2������%���w�,��� �k/}�'��RԈ� Ʊi���`1�i� Y�M>�1g��.w��߰�TlJ�Y�%�S>�<�T�lp'��Qtl�ʣİA��6�9�!��2hA��`s��c����d.X���	�|R5�@������n�o�MZ,j�'I�����pz:�9uf��ũ+�s=��1}��	Z� &4�zӍB�Zp*��5�k)�Ӱ�+x�ΐb2j=�\F�u�m[������FAg�gd~.%���;^�A*�Ms�9(:ī1j.z�����_G� %�2 1sisfoQ	3*0�Hw��	'E�˙�yyMI��+K9DT�R�t�{���S��}�{��T/�Z�A���]B�ֳ��p}���<�kӴ,(3����m\�A ��J�����S����ԁ@��p���g�?ϤZ0b&95m����a�̉t�KA�J]GE���(Z�82�R�S ��墜��!E�%6���hG�S��}y��͚�߭�F�&���e"�ʟ�M�t��>��v��.���4����M(���9C��Sp����Īp>�{K�PR
ղc���D )����>�"n.פk�:тLXwtF���2�Ƌ�AA�1��s����sY	"���`�J7N:x�](6:��+�k�ْ���(��d��)T��l����+`Z+>���l�{���*\�5 ���C��nTy��(v����Fth�f���e���^���~�F�����!,E����jA{�~d.��ǴJE;9Ύ"Luζl��8в3���L)��G'=��^)�a�ש s`�&�Ti�\f3(����֊��T��Wk���ip;�5;���S�C	�¤�=�S~P�C��Y �b���O��9�|�Xyoߒ���������:CB�q$�}n�eH�~�[!i��*|RER~O5�r�)�����O�kk##���W�sh��u{cv���lN/@Ӑ���z;C�R�u+B3ِ~�t�p'QG�#x��M���J��?k��왢#��9d���عd{�I�@Wr���=_2��ĆZ9�ۀ�r]O�����y��>�Ti����*��b���[��U1N�]�쁵m ��{������=�)�	�'~��k����S`���3�Lɸ���	~]�|WB�~�|�~�d0;,�VFVJj#$I�QQ�4�¹�1Jr���eI4��rr#d�Y�WE\��<���I�.{ �&���jf���5��.ϕ%X�NY�=�R�7gW�e׏<�\#����τ���n�<vEv�ڵJ� Q�i0���V��yfԻ,��l��_�}�	�4Gr�bN)A!�3[��sR��ы-������T�e1�S�=8�Q�{��xN8�xM�v�cdl@�Y���AM�(Ð�jyZ�U�i.��+�L�I���=J�"��1u��\�ͩ�sׂ�ǁ��`��?H�Q�S�ڔ�'�����i�&t�S��?ȁ�\`����>L�h����sh�e��,���� ���Ѷ;��p�r4O|o���!�v�r#��	�6_����V��rx1=DXA���Z�Ċ����ԡ���@Y_�f�u!_i�%�b^?�Z��Q�s��^]�X�έ�W.\[<f���-ʖmׇ��^����Pp�Z�u#ݐ����ń4��%]q��ah`+��	/]ބ�Q>b�jL�+$F���6�� @傸��,Zd^9�������c�#;�E���Be�tEv+잫v��	�f�Ϝ-��,Cá�ռǑT�;X4�T���֞K�Oɺ/�U뎃B�}���:Ѕ��dG��Fp⠏6
�
.zT)U�������!}��{�7��o��]�IC*'����泚xs߫|��Ƙ���%�:�Jy�t�����U��^:�򘄼�3�'>a�/|0;�'�O[Ń���mM�[r���s �[%�%�ŭ�1J�dp`�t*ؿ��wk��1���-2<�騞1���zL�ҽ����ݠ�9D�nz�q���H�G@j*�,;�f4hv�s�D���}٧�aͱ��.G�C�@�?�4/��9,�+��3���$����<�j��W���^��n��zW�{$���b��y!	��!�?!'2�cƨm�6k��@����������w��N�=Ji`9�6��ϥ�5 ��7�'BV��M*�V�AJ��ߥL 64Q�a!~��ӢWT=
j�+�8:ϛ���@lE�0��%\����HmX���Zy�_x�d���O��],[��^F��s���k{p�]��;x�v�<�a�6a)��J��"�DG,H-�}������W�^��T��G�k�4��:�8#y�2�,)��:֧�E(��hg�3D_x�Yᴸ�7�=}pr�-��zS��z�L��*/�jN���Һ�m��>��1���0�.�����m~^ֵɻ���v!�K�!��(����(�=?hz��j���Hx�����R����"�2X�`LN�)鐭M�Q�L���#@feiN����$_ޑ%_im�ge���*��u�F�Xt��[!^�/>�s8��Om8����Qo�"��k@��(i� ���k���aQo���Fg`��iQ$h�dQh�)�1��v{�kp^ߙ%��!
cl��|�D���S[�>�}Y��>l��V�h(�'o�ɪ`_o�|5f�6��Ě�g���m'��4�$0rd?�rݹW@x�kp��!,��F��2��_�v8�M�b9������	��ڦ�z��O:���Q� c��^����,��8�a��kƾ�xÝ�l,��ّ�
�fD��g8�������дn�!�Qr�+�"����J��6� O�Y�BI��M��_[?>�(�8.O�9��r�߭�U�B�<�	Qo�8U�F̴�T�c�����\�aɪC.�����a� C�T84�3(V��ɔS�a}�hZck�c	�mj��