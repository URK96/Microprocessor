XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C_7�G�� 46�gb�F�X�&�����J���>���������%�o�M"�l�K<�N���V�4�Ӯ�*�ן��Հ�5R8~�Q+�Bq��WC�`��&��ؗeg((��Xd�A���iyC�ת.i(I>+��*�]�y���@V�Ӊl��(���n�ڃ�9k�i�z�މ�F0z�Ȏ'BG=�m���2��?M�z��p���M*}��,�u�lo�"H1�<�1��c���<��-��$k��j>J����;6�U����)JS<��?d��J�=pgHb��� �$e�]��Ey���.kZ����r����sxa+�X�j4�	@/A�bK��X�\-�r}{��]��|eУr1�Q�Q>��.+u�!�=*~��[~��	Z��L�C6첨��
��i4���2F~�r�0��t�mGބ���ف@��Ҡ�S܏D��С# ��V0����u��r���I���&�~�\�|�!�lh�,/�FD���1�^���$�P��j[�7 ��-lj5�7�}���pO5�/�Z��`���L29���%�U�r��:�/�����>j��!����7}�T�����A,����F��o��T��֓�:~����/=�}ܥ۽����*v��\��J/	��F:b�5�S(H��v!Du���UZ߶�E����"��4�>x�25X)�@��4�����Ҵs����#��[<�Z"�.���D8�׆�δ�@��O=�c�沪XlxVHYEB     7e5     330����=K� 7����?$��4�5��?� ������d�q���~ܤ2��V�j��V���x�l�[>#�pd�?+� L�(��+~Tp�Z'O��C-e��#-�P����騣.�����4�T�c��UZ������:C�n�^��Ru�������Jdi\t~w.)岅��1��L�>!������qc����0����a7z5���_��G�x�J�c�.��=Ba�����U.��F�K�ơn���a��Jk��C������N����	�6<?�x���̥lJ6D���u��b��m���)Abʍ�l���K�f��?F\k=�e$���r�����m�e}.�R8͸���>Y,��R�Z�Ti%d"�U&���qy��߱�F�eӪ^�j��{�^�$k�����T��"���T
C'�G��r{��~�����Dm�u���E+���L���Jm�<��{���ЛbWn:�!_�M��LTE*$<X&Rb���C|�	ʊ���f �թ�PG�8�0h��Q�w<�|P'2F2���uDݮ�<�!��KRjq���-=�[RD�(v2QQ �m0�EY�S�A�Ad��;�:��OC���E��L�J��o:��T���<u�E_�V6*+Ur�e|j$_G.�-"�ᡉ�e�`�x�+>��WU��d'�I����B��}b�C������۲>e�9�s��u��.����2XYݦ���d?Q��Y��nm��`�<��!�3VЗ�..$~P�ϤҙֆY�F���8DQ���