XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��O�h�*d��B��G��gpQb~Ū ǌ%T�����}n� �v�����GF.��Ȅtā�1��W��E'�b�='i�<�1&�����x�P�;�7r�+)�F9q1p�W�檳%�̩n�<�����uu���y5��.=j�zΖ�ľ��g&��n"�+m�@��3Z�"O�������.���#�(��4��Rd�O[f�
��~�#��}8i�i����]1(��f�վt)����t���/�q4��M<s���2'�p���h6v1t+�=��3�J���zSK�$�0�\ӿ����ӹw:]xReoo�DsC}*Fq�݆�e '"�N�xt��m�oq�_Θ��T�����ܫ�s�W
��T"�rL���Y�8�vT��Ȓ�i���y��A�
\��	�\˵��0��_�3��5��,��#c��@�g�F��?����	i�xX���N�wc��gygtSwo�X/ӿ�%�!���J�b���)*��3��o����@���.���"K��5)���ʦV�2N��,���P��~���SDj� �w�.=jӆŭ�
�l�H�e��b[�)�i)�;oS���^��|Ɇ��x(����-\�4�?3��J\��3�_��yN�	�$fM���i�.(�ְ��c��w}p��ͧ�&[�p�x�r�y��}�e��q�i��L�
�5_��U�Y��|eR�mZٚ������9�J��F+���K��n�?"=���F7C������B�s�^7�zx҂tXlxVHYEB    a354    1890ה�zq�7$��3J�`Yբ��a� @��z�i] I�#s��?=�.�|]p�.ZU�E%�YL5���V�.xUSn�5�1pc� ����w��L]���h�޷��`�ZI ��s�ԥ��M�D}�@�yQ=x�܍�Ğ��⻛K)��,M�JE�ƌ��?��3KT��#��T��׆��P*�3��֝s�\�'3��pT��CWO�@�<�]�Y�)V�.':����1J�"�f�-	�]�,Q|f�>�z�iN��!�n�D�6y�a�����Fފը��'u*<p�����I�������GԹ�\ y7�i8�2���"C$#�_k5𰕸�"/uggs��uH��.�Ч�cT�D=b�覥:�a%;�d��ns�T��5�����Ҝ@�-)�y�f�ĳ���#�)b��J������L*ڐ�hu&�Ő�%r��W`c��h����'*�fm��ί$�V������U��-�$R�2*%����UT��9�Y��5��o���^q/C���~��|��ײ��;����P�@�n*_�;�:t������Ό8K������G�c�rY�*uD�^��nK��	���L0|�x�`j�OV���V�l ���C�ʱ��<�5�T/��E]^��h ����Bᴸ��֦p�%��;:��}v�(S���-�S�"�n��IH�9�,+�x�#������$^�SLH���s��)��5K�><Prj���{��#�P��Pf�᭨�f}�Sjhˏ����Я6d�e��8&�Gȹ·iΑ*X�����:�+�3QP��cY��ߔ��^fN�X��N"�,�O��]cuV�@$:�#v��H����M|��ɉ�
������]�-h�W��N�w�pd���"]~����؋DӲ�ɳ?��_����M����F�_S�6����e�8�H����;F��:�x��50~ui�-%o����o����C��{���C��e=�����+���� I��sjĘ�I�H���P��~:�{ۣ��}�@%�?��c{�C��s���|��.�W��Q2�b��;jv����T�>�kmi��(O��������m���c9�W���/;8I=�7�	���U���%iIƕ�߽3��VD�.�}� ��NA�(�!��7;Ԣ�$�M�|�W�����t��Y���@�JB̢��i�����<��N�|[v3���)�2,j�T���nU����$%Wj��N(�3@���jE��H�c�N=���#����F	=P�����y<��^������k1R�ר	���7&�E�+N�y��/�'l_KH@$w���\��qe��}Zy$)Q�E�
*�t �{���Yc�?#x������I�5J��@;���y���NMl�=��⼧�)�~�
�,��������3t�7��g�|'t���^�r02�#)�3��A� ��:1Bl�K����EVN�Z�#�Zzgy�R���lj���.h���f�$cl0{��Y�A=�8�V��ڔJN`�W@;�8��t=zb��v̋���	��f��&�rD�N���:[�[�2�*���m�6q�!��z&���%=4\�H� ��Te�BK�(��,-*+OD(^�_��]Ok� n�A.,�,����������C��F���BLl�GD���
r�s�B�ı��+��[`f[�L�'$C�ġ�WI!���R�����i M�]� �"X��oȃzQ1b~ܿ7�<��=�,�K�#0��ʔ����Z�Aݔ�{�Oi1GO�n{ZVq�ngo6*&��ա�zyd�e��Q#:xoV��<a�n�urV����;���
�ڣW4�G�92�U��ݱ��֔b���"z8j�Y�W�J8m�~��QVg9��+����֛�U�3Y�C�u�D���s�N����\D5��h/@�Ya�e�P�'ʋe�5����~�Cn_:'��H��6Ig�M�? ~%e��ϛ��Vh~�4��[.5_��+�v�#z*�ԽG�@�n��n�8Y�E]�m�:S�!; 8�Cl�Ê�C�LЩ�0&�0���]�Xǵ3`?G%����S��P:k�j���k�v���u��`��8�ao���W~�\�%��*��R��d�%��(�&Lg1��1�G��
��X&��|�d��d��#\>���vh�A5�5�rf��B=�}%����%�7�
�����)�S&�����~��P��*�w9C���+��}R_1Ƚ	�l`��ʈ_����!&��Մ�e�<(cm���?3�l�r�Դ�ne`�@O��U�ϲ ����O�PT�nO�4�P:��0�hPK1D�<��\���,��R�6��ӿ�?��3�̹�NKQ�L�F��́d���<���+�h7%+�S4R�"F!c�����5�c����V^��'=���3���U�V�R�3t�����Yw��l�������fG��2��";(;�����^6�-v-�IeC�O�_�*����fI
%tm��@�P�Ǆ�~ℛ����`�?�[۰Au�
�͛�]Z�4�e@��)&m���׍A#)�gD%�� ^�;�j��+���g�����S�kƐzX^-OB`AD2<.�<�5M�H��W�fyv����0���>��)�}?�@^Z�ࣈv��f�Q<�/TE�$̒�ڬ&���αc:������{)%���R
l$?p�篏��[�AAǇh9M=��<���`:rf�3���݁A�=� ��iJ�},'�tnP�lp:O@��\����A�������5���Q�6��^�7��@9�jcXF�ܢ`�3���(^�F��]�U��~8�8�lY��=[ϼ7�ۖ�Γ�]�̯�A����'�;���)�$bȤ���G�J�I���:p�������m�;�sLL�z�l��X���B��e�;����Olf�����F�[��~n��2\-�k��G�ҔE����'�e�1�g
�r��C�7�7���<��d�*�)OKHry�.+LEچ}�a�	P>�+���&Ǚ�_��ee��v���2p�d؉�&��	)�k�s�MaG�~�:\�<C��bW`�iȩ���}�[�]ĸu�G>�4Y��o�עӲw4��=��D�G�jnJ��]�L9�cjVm{πz�ց�80�lM	p�]��r'�ݹ�Eg�$Lpw���ރQPF�\,Yb�8^W�.4�+H���,���v�&' �[�3���P�SG_l�'���8�L!Z���C��`]P%0{���O�o����(n��d���"�o*��G}=���2vc���n^[���v�ʹy�,i��q���j�4!��@�a� �WI�����.�S���~�`Pt���&P�g���چ��F7oc�u�|E�3�#����1bU�e���=���o��J��0����z�K)8��`y��T��O��p��ۺzM���`�=��,�o8q�칏0����	�o����4����/����_��W�k~�WQt6[pm�����h���/bn�����z@��YbЦ��.������/���N��ɔ�9fG[ަ 	��^aM�zk��!�X=FX ¥�7D�.�6�}�~�3�x3�GL[��d�K�ǡ�wF/04j]|ǩ@�){9�c�L���I>8���iX��5-������=\��D���n������Z] ���^����k�]��]$��g�.��MӢ\-����ڱ?-x.�!����0��Q���K�/�~�ݕ�ݖ�B�(9δ�
߇��ȡ�K,]��wL�Je��'�?�������H}˕v�b1hB�<���f�x�E�������I]�q�2����>�8Gh'��>����Ja�j��Ÿ hT��޵3z�3Z�޲��1�El8A�`����{�E�^E�5��1�*8�(���[e�f���V�V��N��c��~��=�/5�]�ӎ�*EM� f�h*v����0/l:N݈k���%����v�����/�c���^�9U�A�\]~�9��'&>�I���c�����ң����~ ��`�k�	��I԰5��r��-��k�d��NFʄ�mmu�tbش(�h6�k��4WtGH3eY�1�e�/�[�=��Nݷo����;Veg+�#�#/��⥝�aarͤ�9a廒�( b���5DZ�t�!C��4���ĩ�:#3-?אE�ã�/.tlONΤ�5yX�{�6{ύ�[�El�֘������E���V��]�U˳�Wd<��N#r��+Y�(�_BH/'=xf^�@C���G��1Zu�W�{��5��4���@ȡ, �N�19��,J4z!� ���j�����0�qĭ�w¢%�����E�:�J賔:6�,b�e�V�4�,�$������YɆ3�(
*��N���}��(�"�j@�� X��4�oR�J10ٶ���"(
�i�Z��=��c��`��mZ�gn�t�_^�d��818�����3�^;;?2�;,	0�;|k&��uhZ���y@��C�!'۽-ӷ���󴑼�W%% V$
;�3�eu��<��[�U��/�8הBt4u�qgѹp��s���t��a������COm���:��F�p�[�#D�=��U�}���� ��j���z�-Fp'[O����3�!b�A�@�06���"��[7%�	���t���vW@���83��"}�K��flb0(H����+�k��ߍ��}
?���y�\/��ʨay�{w�2�e�J�T�3��w8�V��c}�x���?�&�G����\�Ļ�8���6`O�AU�i�5�����7�P:�|���U��s�A;RTֱm!(�������(�Q��hǛ(��,AWo�F2�0K���>o�2��L����gA4���*�Lt��F�C�1h�\~��5T������D?5��i�3Q�?ݞ��C7��V�ߘ�eO�Ҭs��v��|&�,W�r���AniU�����*�_*��@�3��<��-�l{�>X����^��:``L��I	������W3�������Ya~�dJң��U(6�X[3�ɔ����CN�3T��U��J�R����>�6��
MНː8���%Ѱ���ha�nE��s��xbR`�������;q�ͥ?4�ҋ�~���t��@[�¸"Y��Rw^�'���
�t�P5B��n��ؼ�%:��m1B�#��^��2s�J[�6�5�X)���I�d�k��r��dP��:��أp�㈞rՑ���?��B�H�K����3mlh"�/�R��{މs������\h|���-1�_�z_��`�늝����ڟY�Y��B�Ω����g<\�5���-T����v���x������ؚ-���`�%�mHhX^�5�?��nƌ{����r?p��N{^�i��>�.�Ô�lJ�*qf������خ�X�v��r�KQ�$۱��4�����:+�P����q��Q��ȟ�v}*����ч�+t���Wȓ�ҿ=	�h�l���E׊�0�`��^蓨��x���ط�����I�~`��e��ׂp�����5tC�R��oydx���!/��]J�*.�?����m'&.㤫��\O\f������/W�������7fMF�?��}� (�����[rIR�kKc��+3�ʳ�)�@�Ƴ=����/��M�yÄ�m��>M{iI||p����qq,E|�'��n�����lC�8�p��Ӓ��Ajd��f6���=�-�n���;���8��;� o�&��ݵb���?ε����b3/?�>n}��(O���������S�&D���jZ��D��p�_>E^�虞���`(<�M~�� �e$�{"a\�������Yh'<�k��3h#f�Ew���~�N
U�_Ő�jg��'b���>P�����*`h�H�c��h�y���ߏe���pd��L��辣��y����7�?$'+(��c`��Q~q��N��]���׸�+bsF������t�v�*'+�M�k�ף��e<��&�Ζ��QL��)��`7�X���݄��-�[���ɴ����Z��{p�\���Uʆ�v��eS��OFS'+�Xg�m���v���@@�f�J���惑H��Q	T��}���u<����^1�i��_W?Ġ'-[����i���d�E�AH��{W�	��X���h���b�� �