XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Z�t��Aa�Ep��H*�},-�0�v�Y����H
x?�P�b;D��03:Ϗ�ƎygZc�?r�������<�K
��*0��d>���N�~���xEo��g�Ё��[�[���o2D�q�w�7>����$I��ոe����*��f��� ���vD8z+�đzU��PD*!�2`���a R_�\�[&��Rc����7rwTr�1./@�jI���Zb?f�݂��9UW}���َ����F���������b�>���򌬦A�̙oo"0�sjdܤPqԕ�ǈ�q�-tt��nj�upH�p|h�Ӟ+����>X��NJYZ6\�9��>=d�2	֪�V�V��b�W#�/d�K������z���p�{�.0�V9E��A��5!��T�|�y�4<	Dl-�-O�(��4-"�g!a+��zH�)�fP��L���-Mo���V�SN*V7Y��֯�u��|��%�+t�`$�z�M?.��w��%�U����z��f�h!��.j�}xCA�̬n~��U�_����^��UAC�q!�Hؠ����*g �0w&�Ť8
��4�_M&�;~�L���V�IÔ��g�х��>w�d*�aP�&��r�ܲN<b��������9�(�Q��\b6#i+1(U�����#d#��8b�i�-d�T�w���$��	���ބM�ZrRܓ�\�]���a;�Z\]��I�[ϣ}�dD�K�ͥ�cFa]nD�/+��g-VZ�vH����e�8�ޒ�XlxVHYEB    41be     c40���<��xBn��PwM��-9zM9<$Go� D餖��b=�S։*�G"D��Z� ��78A9��^7�J��9��4�F�ؘ��y��Y-(�%m�l�.(Ue��I5M��(IQ3�x��g�Amw�� 
h?��0O�PRrS˾~\�����܅4����d��R=�E�z�$|�̆t��~|}�c%r���MmX5b�09r*3{j�v��b�	���X�)Cx����W�T�K�+����M7x�z��7�M���{� c�m5�a `v9��ML��Ǹ��mOfE�ȁqǜ�K�yPj�~L�)�(��(<��(��N5�z�s�'ճ��Q1l�d�9dW-�	������.t�k[L�:C5Y<?�����Xs1���@h��ǭ��9(���!�"�+���QSX�.?��̇b)�[: �O"v��9��Up`�_*���no7��u[�
;\����ӻ$u��O�L~��
�����:��/�����e�؜��E:�^�lS<})����JV+�iB�gV�C7v>�ׄ�w��,�XE��[{�b��o��ꜻ��`�n��	�Q�_��}+\!X:WP�cVu�C�i^W��3�{c�e��W�ϕ�5�\O��+?*�����(��g���k�V�0iY�����C[���㎏T�ʗp:��L�����@�/$@VD/���$	XĻy�}^����ҴoL̖iyRV\?|��[�@ r�t{P��R��:���N��O�k�o�����e��V�s�ߤ��Rկ���Z�1�L�lr���u���vo@�#뗷��8xÐ������kV�^U����ȇ��Ò萗e���R_��>t��4��w�RP�Q��'0�]J[z�*LN��vdkƘ%�Y���H�'Q+�9����$��X 0|���g��t� �^������o7��`'�U�HX��a������r>S�}��
AK O_��(9h �����U�L�mu������� `^H�_�mrx^������f
h���]�z��⥪��#eC`m�O���=+�����u(�ā2|I8��x��kroi������ja>��9(适!E���T�(glQ�3�}cX|�EH�9\	W�~��L&G�ѭu�+���@�xj�ëe悆r������03�MX��A�~+��S�r��'�N����˥�B��Y��+���P�����wN/�g	]bHGd��I{����@�?De���*v��J��m��1�%��w3�(�j��'����u��؂h1}����Z^�Pq�"
5��,MQ�:�(GJ�n����Pmgz�������H��-�_\�I��9k��М����Y>,;�E�f��%@��o\N����A���v�+���Ag���tx�m�Y�/B�l+}L�Z�΍�y�X��$bTq�l�E��! ���d���"޼9�ߺ�@2%����"��ɰ���~u�i�>�.���.�㗻����&������0�L<���3՜����К_�,��h�%��a�Mp-��/���D�wL���4B$��NJ�p����˝}v=�榬�֐��/���7�Ff	.��Rsoad��L�bD9�K�$3��Y�vE���Q�9f8h����k-<�ְ�)����=��@!��¯��1�W�{a��O!,0����m?i�!�ǎ��,76�:�АIU�F�J	 �P�f�S|���'�%��R���SUM�1���w���%�q� K���A���k��q�Z� �\۲��D~Ԩb.^�+1.�lQ��j��U����Ŏ	UhE|��D냗k?y�rW����bV5�Bs����u�u��6JZ�w�, ��f0Gq0��]�?��K���x��*yU4Z��8�fx��n��*�5}���I/��X�%d0�!��#�x���r�J������)����7����?l�C���}B�_D�<�'V52;� ����¾���(]QYΉ�d��Up̼-�J]���_òxĴA�+��:$�~�� ;�P�:��*s6wHf:��\�^Y�vE,��g�w�C�K��'S�[*��?tz��B����=^x!�����s���n0�M�Ɍ�+�jG�9����t�!Da0����vE/7�H ��s���3.�dk彁,���vr�����0�yWm��/a �M�Ԝh|2]({�Hz�:�O��3���F�ٚ����b{;��#O�� {{��H{�����������Y\'XfT��6�~!b"��z1���
F��_�rx�H�̗>��l������?0��H����sG��1���"8�doA_��~��uG�>@�u^Ko������9�~&3���xSDo�a�j�L�f�v�A&7S"ˀ�`�>�V��;���?�=6۫TU[�b��J7�"����܌Q�_�g@i6�_� ѵ ��y��[��D�՝����+�%� ~S��0�(�x����0Y ���8�3 �P*)��
��c��\�ǆ�-2*��3�D6Õ����~�P�]�ڭ1�lGD�	�ƌ�F՗�����8�\R��è���${ք����13�d뢤���-9S@����Wq_ �����8&�#`�tt3��uIOi,RV&������'$����;�F�g-�F�;�3XJ�5t��o�$KA�!�H(&r4P��T�ئO�m),:��f���8B��3F���\�!XZ�'1?Ѐ/"���F����ТN�A��8q!g��|ڤ�n�0"��/���[O�%y)�Ki����R�ic�σ�w�*���A㛊f%���3�֯���T
JR=��|'�f�Y�y�<��ZhO����i������g~ ;]��'�?�,�JQ��T?@�u@Iј"<sha�u��k�&Kr��� �@�+z��K�>�
�\s��#hbh<��YJ<��~`(P�����,�#N�G�IT��n$&s��Z�yٻ�����T(��<��Jo��hGC���>�C�־�.�m��o-�K��� ��ѧ��^�	�	E���Pp("��(������w�1wx��Ӆ���-L�.�U�
=�_b����i�}z>iO��S�ŗ!�{�%jDы�E�ds���