XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\MU�E�{�#�q�TT��u� ��ArOn�Y��溼�eߗY��5bS�1�X�[�k��%uZig��\���ݡ>��+�So�Y�ӻ��YP�4��	���.&���h����6�,�FbI2J�+$��E�&f��T�ء߄���e������)@'��Y��3Q��!	&���;u�Tb�7�F���pθzo��F҉�F��R�S�s���ݻ�%b轘��*9 �hc�����[V0������7�WJ�J7�1a~r�o��P�o�ê0m���7� ��doy�D*��9�UU��騉x������ �܃}U,q�o����t��C�@�%�kV��eW�41�<�\���K��Yp�'ԓc����2�,���z�����4'U��Vۈ��n���=�J�8�W�p"`w�4�ds���~�k�c�=víF'���#�~pb���;[��n��-I��F$�a?�����ӊB��S�������>^�	XS�u|��v	�1(j��������.�3?J4!�@�Ϭ2�3g��5�~ �6_NK|E�>����#�z�1QO���.����the�'9����9zw�ޮ��I#X����� �i��o|����ڷB�<9��u�I��?�|)�R+Z ����a�t��@#��0�Pբ���(�l�@l�f]��%��P�.�F�[��xE[`Le���l�tD�)��E
��M�S��͔���h��qF�G�8����XlxVHYEB    1f8a     780+���kSE���5rSp����K�a��]��+ ;����B�wF�g�1Y���H0DjP�'ڠ��\1U����m�cy�����`�pDo�\�Bϕ�y+<�>�)<=NMxM9�fT�Ն�������Ȟ|��^�f�o<1����m+�
.�u7�C���`m��Tr�^����0�J�GH�����H�� *���<+Qj�����/9� <ib!`&�������V��IV�z:_�g�9	�t1O�o�L�C�`
����er/��!,M�v�c'�U��>q���Ŋr��1	��Z��B*C�rTKq��X��� �P� ��2ߎ�X{l&�g�d��$}&쿬{\I��/�fYb�x�j���^~�ZT�1B��M�sQb0[tg�̡)�ڢG���:�4y����􉋊]6�e,z�P5�;�T��Nko�`���t���v�"�p�L�]�k���h+�:L��h��^z4��m5�43�(�C��AG2���Lb�A��cT�;[#�����x��0�Y&S:�jQf�y�}������_Z`��Z��� *��ܩ{��W�Mi�.�Ym�4��s�;��!�:�54�c�	��!�#	����!'H��)�>�y���#J���;����aC�D�e-Z���@ڗ��uL��FBF�D��y��
eo)'��^[ZsUyϫ��l�v���i	�k��$�u�:��zɃA�W~l�9
��[B�ך �v_���p�"='@_l$}����,!3���_����0��Ȑ��no�B�&4��q��L�A�V�l[�J��~kk�k9B��DW��L�_,	6��4�.�1��枫�CL�u�f���O���d�ݛ��
'.��'��FF�ȉ���,��_ �a������8%o���4�1��|o~7�T).Mk��c���P7U��	�̚R��HyXש��BG ^����N5�044Bl��V�e�c��� /i>>�b�G[�%���Q<��,s��V��%�@�>ccN&�7�z��:`� �*̑Uβd��l(�-ZA|��B�?��$i��V%�:6�����8V&����EN�����(. \g4����4�pfc���Fb���m��Բx0'�x�iKZ���8B=/2�-�1��y�2)�>,��(x��,����6��/�V����4{vE;�[BY�ɼ( �<���N���A�}��x�."2�o����b�-�7�Z{ۙB�Em^��z�ͷ����$%�+m�m��5
�m��,�{ƽ���݉6:ϫּ|�V�:��(Џ��5�%Y�/��_����}������c1��N�z�~!���v��{U��ꑆ���G	���p*�]m�, <s8�����4n�ң������!Y���Y��6�fw��	Mݫy	Rxg7��46�~S�����-FF��6:j��	������7�rV�B�ù[0^�ј!�*#��_�=bԅLG��Y��Sp��q�9�Ӻ6h֖���L��pnƾC�A��,�-��V%+�ЉZ�&������^�.��,@��!  �x!�{�c��'�(mM��r��\��]l_D�c�z�ӎ���"�ΏJQCJy[A����3�R1����<:G��U�4�'�!qJ9�>�H���/���˪��LI�mx�C�U���_q �T��ؖBh���$'��2Q�Y����a�k�ɝ>j��Zͳd�sBx���6���*��h.�f,¯D�ޭ	�#k��>cPc�F�����C��J�M�r3�q�Gc*pɋ���Ƕ��X�[�fGt�].3_l��s)��ى_���lR�s_ܧ�n!����C�R`������v_�-�C����#�	��#���m��i�