XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��DV"�i�W?\���g��B=�{9 m���j$!�?`�׵�e��kIv���<��vZ'�4�HF[h����GD����I��S5D�锍�I�LS��M�/1���8����31�3N����.l�diA�Ń��C�h�P��D=�Bc�;Ih�D}W�0-n�i�^����݊^�Q�.?� �G:ci�m�g�Q�o)��Hvw���	�W�$��SD\ߌ=aj��c�O,sbwI�[�|L����� 0��G�` 5�%֡H�š���<�R���U��83_ �E�@��i�`ĊUП�
�9Qp�Pi*+1��^��kw��ىL����O���w�D��^�]
ٷ�w���|E����U��Oќ�7�z�⏌�RX�X�ܟK��6����8w=O���%bQH|2��ܙ7:s%��y'%��q��ţ`���=��.��	�٩cs��)-Ϙ�r��k�d}D���[�oD���F��AB����H� �uY�T ��]�ѳ�"����awk-0��Q��bɊBtf�&vX\}ѫ$bz:�O�\�	��)��qV��Å ��i�\~%ep��1���z��_��8_��$4c O��َgG 8���7������0u�h�py�p����x]�6;]���+��{�14� %��Gl9\<1�.~H�����qQ�5%�`6z=2�+��Ҹ+Z`�&�T/���x+'-o��L9 �����,Z)k�@>�	DF�M�S��ԌQ�($N�XlxVHYEB    17a1     680�̶L�W�YwQ=^� $�՗,��I�mfQW��aV/nC}!�44�>|K�-����!)���Y���g�i�pO�&��'�o91�#-*�Wds��H��+�"D�%����R6��_D\FE�C����w���8r����uz10���� h���`r��	�ROO�a��6��rƸE*Zg0H�9����L���A���=sz�E���0���h~��Q%*�陇g;�2�*��O�U�m��5��^	�!���J�F�й?�q��P:��]��AS5��^��ײQ���tT�6�Q/��{Fl�[��9^��jD������z�\>�S|��$��`�\�g�t�OO�:�;��+XSe_+��62�N�O'`����@����M&rw;;�e�_�P>x�2<&K�����x%�h��&�������K�O�U��ud�{CD�e�粐�)����,^�� #$ �ɥyd74P�KA&�~u��C	B�fZ��	�">*�`�D=��Dȋ�'kj�vG��3�ڤ`\�vD|?p, Q�{�.Oʇ�]K��
-x,�Vl����<<f )� ۭ�8��O?�lC�AE��h�5)�>�7Tо�^�ße����I[�w���`Pq"���J �;�Q���4�b��M��t�lҢ�A�y$�jNnGo�ak;P�o�T�Y��u�Mq�,�e���,�V�%�ID�L;C3��W��$l�XA��h�֝�r��4�.���m�vi�<��X�P/A
LAE��������ϭ3��+��]���K|�8͝���u:p����F<��2~�ZsI���)F|���
��۳��k잣�k�
����_|{:'#�k���RZ#/��9���L9�O���2Xڹaݾt��s];�0����(+�t�/�n�n@�����X��>\�BB���0*+K���*l��"�[�2�M�Z*j�h�7�J�yiѠs���G���hQ�!A4>'BR�'hg�e�7�,���b�c�t�0Ȼ2���*�rJY^ƗM� �������Fΰ�vP?b|F�l�e�up�\a|;v ����;�.��z�
/6B%�dW����{��!�*�V (A{b�˂ ��	Wk�.�ft�9��$����4H�k�U�`���Ƣ��c;.����=(q�[4�V�ԋ�wr���R5��3�*�M4�6����d��K��W�^�[��׻vl���HA��{�F�oU�����o��^t�8-���A�d6�P�v�x�	Rnl�D��P'�PY�A��P��i�G�o�nw�����3`�B����Wmt1>�����"���ֹ�Xu۲�_@�Uz+$y���E�E$�%���2���L�7͉�V|x���9���v?����~����O���7Vxl�M�4��o
Jd3��w�J�1�Z�=��[�� 1z�WM7���5�56f�0�����7 �&�3�!�N
=G�>tUC ���
K�?7���	���Yz$���>�ZQ����8�r5�iϼ�|��U��B	w*��J�0��h�:�S&ec[��k�N9(��ė�8�9H>�U�ڬ�Β��윁�#�ӶC�X��Fn]y[�:��4��,�G2!=0�cvUOe����#$��7��v�Y�bm