XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I��E��/j�LpPm�UL�F%��\�z����r1�uF"a�ZAG�z�bF�sVL2xU
����Ǥ�x�C�ks�b���<b:'��<��� ]5QBON�g4��1f��*
u:�M�bM�u�H9X��B�tUF
�K$�P�OD���,КF�l��pV�����݈%���<b�\d�P�8���o�����y֭���W�!�[�}*��9;�(0nɕc~B:�r �;{i�1b�`�"L���0�c��ј�Vփ�T��Px��P��f^�����ZjO�xA��:<�Ė:>2T#�q���K�TU���)wʓ�GF���:K���w�?Щsf騒�f�o������j`+A(�9����񚺀;��E�tdnS���]�T�!�o��7�;��d�g��wRNז���g4�*���F����A��,����%aq�٬�V8��ٷ��t#������P�"cKb �iw��D��'��s����LO@ʒ��	���c��g�6���u9Vk�͌ٳ����B���0���d��E�g5������bky7g�P���F7�4�����y��^X��
��y�V[-1�q7�q�(7֟<8�|\פ��^ox��UZA�x�J魵����WL���=*'�΃�6������N<�t��W�L�ެrw��o��!ʭh(#.�D`�i���<��Z�](R\�j]���o�R�`؀��D�����bS��EW�`d>��m崙���3��XlxVHYEB    1902     7307'�RӼ��J�!ѽXduV���'H�j�ES�] ?j��%��g�[� �t�����A٫��!����'W�Ea:��h��u�N%V��1�6[:ϋ� �H������P�I���B��ri���/�	S�5���˟�9#A��t������'��F6�@`�1�OsE�bQ01��]	�ځ&#�I���.:lȟ0H���G5��CغyO=�S�sǹȌ��v��|_f�ȤC%�0��<�/�D� �(@���hA`�~@�Ȝb7q�������ʩr�=�V<�a�lK�	����5ϯ�Zf��`E�m2�8���S�DQXd]��V���n ���x��z�uW�WQ5y��x�}�>�-�LBq�9wjG�h����7�I?GZA�!G�^��Kt����Q<�bFQD���[������`����Q�_��{�+<m*���a�5�C�e8M.(�zs�J;��JDω�)��bqA�3�}@`,8�#�0�+խ�͖�_3u�
5����Ng"�0��J����ί�ѫ������LN�Xz�*�˕m��;Ĩ�0^TMM��f������ߝ��F�4��=�JЉ�B�q�<b<�L��[5�6̘�,�YuP��d�Q��>�!\imc���,�6�wBp?{��6�����H���+e�k��z#�%0~�T������zO��(�QLQ���j���[��\�P���)Rd�eg�u����ԃ�Ys�L��4!����p�/�m�*����xCR*k;��lZ���h�U��a���Y0=B8��4G�s>�b�'7�q���zޔ�������҉�(��N��]!4M��$�c���6)��q�p�Lۅc�=E��9>���X�
�r������q�h�񡚕�ص5��:� ��$��]}%	�+�R��;��`�5Q`Y�1�f�m�Щ��Fϫz�)q�H�
�~�t�Oy^C���W�q,6#G��k?8 �ϴ��R}�4�Ө\�U���Г����G
ૌ@���/ݧq&���2���"��i��W�XfϢ �Z}�AG��а�΋����a��J�h靼�!�î��WY�f�{��ge�{�y�S����)�G#K�Rbfq|�i���%��7X:��V+u����1ZiP@Lk�'d���� ��~����OFG-R Ɔ���|�ɥ�M؆jx�P+�bJ0a��5�� 9Uƿ>�%[g�*q�)����%�U����c?T����Z�0�u���1���܍z�����|�����&�3���{�}:����vԊf����GA�C��o���caE��(g`V.Ske�y��J�J��2m�ڏ��!�Dw���@�Ĕ�ǂ�}ٻ�IxA�����Y=T_��7�
���/G�H{��@�q���'�6�z��X��)��=*��m�Kkshl_|�;�R6W�z��Ϊ��p>ڶԢi(RC��e#!F�s�V,��l���b�(R�T$t�#j�����3U�H4���pڣA���5�G)���:"��͗t��r��X�R7��y�<�oW��ݫ�`���>F�\�Iyr�Q��/��,�����&WH��Z|���$�l�����N�.Q�𢐉��N8g�pM�]�e��L�&O�}|W���s�i�<Z�$�%��p���j����ۿ�.�8f���&N���x{�*��2g���Wuo��m��5&��O\q���9���-��8�������-f�:��u6�/�̤C�J2Ut7WI��s]%�9���Nnx��@Qif�����R;�ǲ��C�J�����h�qO�y�n