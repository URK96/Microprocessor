XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���r�dB�B[�!P�\Ys�{�3cRn��k���Wt�I��t���$x�M+\L`7�j����
��f1����k9�K�	�����.�G>lw�E�J���sh"��ϑ���%U�Ķjit�]M@�9����_}N"i�$Gό,w'��W��c��Ы�h�m��������$!1<�L����!���ڄ}����U���Rc��S1D'���<�{]������030�jƍ���j4�5���c9v,9�;;>,f���ւصj�n�gtC������:�X���Jߨ�2�g�@m̟*�AML,u�[DQ�%u#�,o�.��	����Q	�KYi*��h	�X��hΒ"�9hLP��P�~F�A�L
��!���[�-�!lr�}��d'�2(Uۿ�Δ9WZY�{hM�[`6��PA'_��b-��ʔ觿��>J?��	iX�i,��W�X���vGDʚҴ�L�I�Ȅ4��3�ҹz0O�YTV�c�F�n
�� ��9�!�[IB��,�d�:}�l�<�H��%�95�*��<KlE7��ͩ(��d3�%3�4�6W����;�J�L[��ݭO���r�c?�z@�J3�E�&U�-Iَ�lm-�/`����dh:���-��M����z���? �O��]�Bc
N�YVV�=j|#� �M�"7C<��h{�@mȋF>���l]��r���[ 0G�z���$���~� Ec��Ij�LI:CXlxVHYEB     7b8     2a02�(���X(Ę*2�l����#�捍���
���ʘ�$��K��7l�l^"�g� cd��m�z�G��U���J3G*7�q�J��$���^���2�fX��=ٲ>5��ҋ�	����V#�u�g����*���n�>t�%���_���IF`<����w�4�'���xk��L��3*��쑞Dv��
�߻q*��;���N	�ݖP���y
-����V�l��u.R�~��a�l��aN䷥�d;�;3N�7�V�0^M#&�	(�ÓV]�Ju��*�s��t�\�3�u�Ճ� ~�>}�K�V�x�T&ʸ���*D;m�R������E���ʣ���;Lc���j�'K���k��|��?V��`E��55�3�0�UXb$����x�� �
����t<�Ӽ7�RsAn�"wm��rb��e��Qf���,�� ���?��țf�0��,��2�}��O뾸�ס��� ��:�S�}Z7Ȃ����f}o�|��
Fz�>�wU��:�Y���`��)��*��c�y�]�����ak�\I��%����B3K��g�f���i�T��'-���i��AY�VG寃��(��|��`��z�q�d�w�_�ٮE�?.аw"���L!ˮ�гb1�ѣ��=���ln�r1-�n��<%����
ok�7�