XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����(	�2���`��V��f�椇�����1ʅ�m������gc�Q¯j�)��}O>���U]��_
�q(/o�5<��ǨA�D]��B�}��S�c�#��v�d�Y��:\�[�Z/��,�h�8����y���7��T���ʹ�#�W��DM�}<R�C8s4�Qf�э��J"���Jky�� ֔P�C���J��Bc��1%Dڪ�X���K?�A�6<�t+b��I�V8����A�"٘��I���JB��\~��刴������F������v�;��Y���^��-����W���|d5�ak�G�	-?_���%	��ȵ�ז�;��3�oE���n ��.��|�뚡��lz.t~���F�j�q��(�9k���6�P��DJS尃��(^V=|��$d�ӛ%k<���7�
�M���_�7R���Y �����0rǭ��ㅁp�q�ìK�S��hM�B�5r��8�v1�>��\M�	Q���Y��"�lW��d��=ԡ�֞w�����UAM{�"R�u��x��z�V�÷��q�j)l��;L��:��+�-c����{uU��7�-v�
G�R^�i��Sݕ�:n3y�ǎ"�nDZ��Qv�G�p��{�=��~ɦ��IH�􉦕��.�;���#��?����ܸ�?u�k0����7��oY#͂�N��G��\ �� ��7L{�}�uv+�x�<�#�>���o��,	�)ˉ��
&� 2��XlxVHYEB     a3a     370U�x�,���Xp`K��?�a#�@�������vvc��(p��#:T`�\bp�Yd����M�&o�N>?W�ge�����e���
�`bt[��VY	Y��'�8���F�(�~b��V t�7q�s�$X�b��sP�aSγ��i�ڏʃ�lQ���L��0%�BA��	#��8��v��C�*�'q��$���gE�*h���\a�n�����.�$��Q�0�W�Q�KBZb�$��T6Y�K-E�ߺl~�<����|q�<n�Ž�(V&��U����s������_hЁ��i�d"����*_�ZMD����{zŷ�V5@�>��hiR��L`�w��2��Gau�n7����r1�[��7b
+X'�1S
��W�)*��lv���O��AC�w�_�^����!�_2�N����5Ȣ/jvE3��7�_g-�k�yb;��1���MNT�R��$��1����%�3�#= ��l���8k ��a����O��
�)�V7�U���dȉ���5�T��H����u�
��󥽊�֡�_"�@�S��l�	�+��66�u$�z���6��O�J P,#��w%A�gw���ܘP�_&EZh�a�gR���xx��tj��c~�,��mF�59�8e^#��Q)YCd�%�w���ؒ�$��h(��|�9�iQ1��XH�iq���2m�p1���@Y�Vs܇��~4ښ�����ᄄ�.�RV$�/s���Q��z��2�T�Ŷ���xw�XءF����($�I8��u&���`h��Z)a�l=�������M jK ��ٻӀ���1AE[&ʠ�a������#"�k��4]/��'�GzssW)§������2ɅGY+�v�����s3b�����6�