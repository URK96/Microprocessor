XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;�!9dw>�b�t�ы�����x��u�K��-w��X��
0LCk?<���}2'.5���dm�SH��[?t��a]����R�F8�{$��ۂb�����TR�N�1Xp��.~�޼�J��F�D��0w6��G_���ɢ^A��\��s��h�H.�U�B��-;����2�N�ڌ �Ƌ���*&�d���M/����]���~�S� Nf�B�3�J� 7�D����ΰ�6�ei�&-���ԇ��)G"7�ޔG��і�{\��ٴn��	��=E��g9�-�k�E}*��h�QJR&���JP���{Pms'�U�Ɇ�m���5/�(�X>`�;"��9����,�l-���52뀔��/|����L1aí(�(r��m��@f~�E�|OOP�X{}�{~z�_6j�?�ea�H���C�y���J�}١�TH���7���{�F&��_"���5W�/�PJ�nwL#s��z�^��/�nf����e�?�d�\�^��˃�N+a+˯���W�d���jJ�h�*<V �������ql�W-!ׅ��jФ���$-����r4\fy�U鏻�Ǚ� P��PD����i�4+l��x���/����{�sK/-#ᮯʚ���a���i�7ԽMh��~o��7[rm/<P�W��Z��`j�Jt��m�b(���Z��UUU� 'JԄ��#R�h��9o�ޜm���w��E�$)h2
�K����QZ�h���2AcoU�lN�[�Ŋ.Se���j��H�1f:ʐ-��XlxVHYEB    1ee7     570V�)�������͋��I �X �#%�hVIx~[��a����Iᵴ^w/����I+��,�ٰ�Q��x�Νqo��?���'*4�z�:Ljřd!"tЗ"���P��Q���)�z��W+T�;��ԱG�"(,���C��e�B+C��ɰ]��d��dT°�)��"0w�b�E��*�o��u�96�W���kG�q��3���رP`����S�4�f�&ĺ�;_`g�k�P�9�k����z��.�Li�]pF=JA)�E-�(�_8ѕ���p9ݟ�t)�e��zu���������)I68�f�a;p��nO�x�؂]C��i����\�º�oֽNDv�:�`�_A�� �0�[|5-��O��ch�����vw@���+tw�,�u�N(���:,�?b}�X�mJ�Lw�
ɦ�?s�Zk�����`8ZP/p�����]�k��^I3j���&+'���S!�D'�%��:�R�
��1�����E��8	z�(�n��0������XsDuьeͫ��K�:/���� ���M4��dc+�D�F�s�K*��Y��%��.9f�{ؕ9x�e���r����ߛ���q��M\�_��v�d\ȑ���07~�*�~$$S��S�L�ڝ�������'%����2�@��w�w�ڵ�h\��m6Q;�Hm�0���c��mN��^YE��Ǣ��̐�d>�@%�Ʒ���jX�eO$�|+�(�����8��u��O�4������K���35�]|I$�(S���wZ��Vμ0��+JQbo����"�z{a:�eO��X����7�3ƻ�m�EDӏJ����~�����O/���|hD�����f,f��#�V9p����x	���KU՞�b ɹٌy��{�w����+>+�Nc��ڊ)gs	�&�rJq�H�/h�i3�$���9]��J��m����dTq��;��g`���8�z��Mn�%K)-8�3E7�/�w
�:�����:s2؏ P2
*��~(�Eb�Imi���R��Џ
���R-k��w��4�1T=xȑ[r�N�c�s�iҬ��&�.�P����\V���ʯXjx
�%k�L��9�j�� @)�s � ��i�I�u��7�"��X!�A�V'�)��A"���v�㟆�3̠���a���^�a����fuw�;��U;k�]��z�r���	���ӫQ��%[P�d<,C�Wԗ�ŨNS���H�� ��Bk�*J�R���TNx��.���Q��[չ��{T|]��+BA���=�Yq~�E�YM:�C)���+١��4G�X]�'�ix���٤�m|g���X%��nw����=;uӧQjӑ����u�p�J�A