XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ս;�"���[�!�-���F��y?y�4s��
���䟍��b6`�!t9�h��W6�𼊴/�/w?�t�*�m�D.�gw�Eۊ�$&^���N�J�����\�rIÙa�RC��A2BW��N�?�(hV d~�'w�~�"��|�b��I��G��k���������K�.�tT�OX����7%�%@!��;�֋���#��&  �-�m�2�E�t�{�n�{��lRG �:�����'�Y��l^=�e>���e��w1K̑@�:�슞��A�L	�=�?~�y@�Z&;v)����1�.��G��XD�tc��tא����уkr��g��:hrMv)�}1�%���(H��Ei�bK�=�GA0�־=N�W$���7�t6F��9�_�橄�TJxNn��
����ٌ�$#���>){^���'Z-Qфm�ð:r�����?�r^#�.�+�!�Z>5
�h!�[����/Z�j�g�^/ U$��	�"I���[�{?��xh�ot��a3�+��D*Ê0���Y-��I����!cW�Y�QFġ�o�q)��5��t2�*�4D��<��>�o˼d�"E��l��n�w]���2�&�ߏ�\/�z��Mn6~"���Z>���V5�
��n�P�|��t�]�tg����жD�^�w�sE�|ZT�n���� �Ж��=
v��rzu{P^�г�xe���#�'{�N!��Lq��j���S�\Z̑�x͍���cnp�.T��`����XlxVHYEB    88a6     d60(��a�;9���زV"A�/��n+����>魲�L;�i�������M$jY���h��B�8p�9vBj��{Jߛ���w�(3<����.�L�����`D�*�N3T�"_IPH�a�?3~�0B14;X���vO�d?�ٙ��Q�ė�*/��4Ta�I�^�\�i���zva%-;�{g��*ҍ��L��֥K�G�6�s��k��B��r?��� /���Yt	2k������$�%���yp��}<�g��rt4�&�Sz�;b�*jt�����.Ǜ�ȵ,S��<�J��O%�ڎ��kV�Y7��M��FsBh#R��K�Ә�T�yۨ>���V��㘚Ҥ`�KZ ��ft�C��A�LћJ�}O�d���	ޙT{8�qICuQ�V���V ]��u�c���%�+Fє�X���=0L���N�b�"�ъ{��bљ����+ԍ�w�:쇐��3tY0����X1�8�
� %��,d��
��v�%��MV0���k��3�[#�ǉ�:,u �Vș�$�2����b���2q�Ÿ?l��~�`�V�n^ݝ�.o5��s��#��*�4mxf:_V\Dt�y������qKu<_+��B��39$m��8�%D�dmQ��c`���ɣ=�}�դ_fB�6fbpB��{�4�x[�˗t�~�b{W�o/�\/K��m�5.�|,�v��2wJm-�^�3g�b$]�7EQ��يbr_@7�Ǯ簊ٰ�q�,�'�����>�?���r�TI���7z�v0o����6_��D�A��P�:)mq�����c)��2��H�_L�����}���xܸB�����\�#����:OO��g۞q�4ݝ�������:�(�%� ��5�Y�P���.���Zu��xx̔	�"�G�+��MOxK�/��0�;)���q�QAՐ�*���V��'�(��
��>��o��R)�a8�R�L󠸏�7xA�����K2�c�w�|�]����L��/�-��G��RS�S1��l�)@ V�oJ[wh�0&�.,D�m�Ǝ�|�����Ӎ�W8G�b��m��[n�o\7�쐭�� ��:�29:�֥��%�Fa�) 蔐�ѹ�D�=��3�eL}��(�e�Lv�y/`��΋��᷎�\s���/���3fi�42�3Y<�hp[��3���|�)���e�^,F?�m
Wa���	l=;��RP"�G?�1!c�̽[�)B�J�9-;�	�K���S������� ����'��ӐL Q�*�-�2Χ�����2�[�u��=�fą)m���Qʔme�i�'�������3�i��!t����ܺDP��ͤ%r�{��L�N/i��A=�4#'&O�%N����D"^�����)vg)HNm^[trn�`d�q�����XU/���l�����i�7Z:%�o�4�9�/��V��"�g�����9Ɛg���^��[	Q�}� e	E��as7�_+��L�I++d��M�˻|C�%O���!�5V�"7IbM�ɴ��8{	��g�(4?��^����팃�ZF	���	��sN����p^�ǘls5n���#�j�h��q,�K7�D���(��}�93�u-G��&��pꌯ:w4�	0f���r�;�����W'�l"��1����t.)� ��[r�jV�]�W��.B��}&�ԋ�e�lmJTH��^�Q�-��'-7���[�����db٠`��W�S�n$b�.��
���B�EO�tx0,���2�DG�����bÓG�X��� �P:4y_�b���k���H��1�Zd3��.�8�d���YK�{�͍���ehuoi���F��J��j{�燡�;�{�|�l5��u��F�Ρ~�)R�Мj�)�#�Bb�;t�=�����q��a 
�L��v���75R!���W�o�r)&�:\��1D R@���0z*
���V���#c�JcIi	�&M��gz�k(�D4�,n���7����;�x�p��Ct�Q�������	�ܠ»�y���w�+,=�67U֡�w:Z.od	C+��@
^+�>@aF����[O	$���ɗml��
�Nծ���F,1�yG�Zj��];��\i	��}��JY�7�&�/�+M��;�ׇ�)%��3x�7�&)H��&P0T��Ϥ&�/K�.tq��9c�"Iͩl�~]�+�4�P�^Ʃ��������~�KGH�MR�\/���86zڻrgg�jRnx�X����Dܥ]o(u������Ǩ�r�|�&��NY@�8� "B��c>P�+�:3�e���w�*�i>�U�;���z��E��)���j��)����1/���vm*���I�p��ŏZ�VC׹��ؗ�Xx��l�f=���!k���-F�x���!���pj,�WC ���4*�fWbawtj�{��#Ӿ�9Xo�M�'�Ws!��w��]؅�
�%�3
|BU9Yt�r��h7"�L���u:S���,�*?3�m�x�I�5L�Ⱦ��Զ9�S��Re���y�uV��붂�V�S�S� �|���+��m�\p���Ni0��"����(�+�ãF�ﺓ��9�h�����x��w�� �Tc�Ӿ�p�w�V�o |�#'��fa�Y�y{�$�se8�����y���+���Bǭ�5J���x37i��i�H�_�7y1�,*6[�[˸CsKZԡ5�-������f��M9X4<��Zyz�Z	�8�,���kjϮ) 6��vƛ������"9ۅ��cYe�S�oOW�<cђ40P�
�����O���w�h��F�2���%"Si��P�UA��^Z�ov#P=�*e�pdV�n���x�CZ#��Wޘ �p��z���O���ڮ��Ůd��w�!n�u'g��i�`,���ӥ*8��������Ͱ���Ŏ��tF���8�mڽ��v��T�"��#�g�J�(=.���PAa,ܻ`��=Jw���J�Q��ٱ�/�t��{�\�=�Cb�^C�<��/��Fq%YF3f����G4��&O]D��'��$�(c#|'5���˳侂m��߇ �\�saO��
������~�y0Oz=g�f��gdx���s������6\�^�!�QU���8n���f;	�aa1�9fђ���!�QfU��[e�����yW�E��/$⨬�`B�N���`�Ds0���e	������l�}b��g>l�5�)��@��p#%��Mz	�<�h���?R¼�h8���i&�]A�K�c���w���&�Q4G{�QGb� �,%�����,{��$RM�[�vTj,��@=Qќ*�hqel��Ig�\��� �fP���%8G��:t��s̜/�wh/��O��u+ӡ�q�*7F�)~�#�?