`timescale 1ns / 1ps

module RAM(
	input [7:0] Write_data,
	input [3:0] Write_addr,
	input [3:0] Aaddr,
	input [3:0] Baddr,
	input CLK_In,
	input Write_Enable,
	output reg [7:0] OperandA,
	output reg [7:0] OperandB
    );

	

endmodule
