XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���<���OQ]����&���<��g�$��~�zs�r/e�7���%q[���с(k�ӕ(`��'����ܥ�$��v
Y����lO_�`0�X�� *�#-�V�y��'�]�!�|lW��2�<�Vj�%mw�$\��uAKԫ1��ɦ���x[:D �"@f��">swa��m��Ȼ�%N�ޥcO/Zq��	�rf�_*1���c�<��(�3j���p�������J=��ŷ�}.$Z���"�4���&�}YD�8w�+֑���پ���ۉ�p�{
�J%�eP�[��!��L���ԅS���#�n�uYRl�փ|��E
���:`����|�x��$3�).	���=��)��ҩU��NL��>B�o���{s��^+�����$�e'W�i����:����+vYn���A�v������鰆l#��U��YR���o[��R?'�H��j(�V�X�%>>���?��J����GxiX���3�	�.:��E�
����ˢ�I�+� ��X�s�/���� ��׬�Wa��k����{4ҴZgc���'"�׋�5��&�n�G7E$�R�����(�B�'8�q.�&'%�Iâ'�.�v��fKQɬ�0�����N���W��AîQ֯��e�3�V���m���DR�uk����צ��ӑ
�~Ua�+UR-��o��-r�n�c^�@%<�e���>٠��4�P�xm�Vߪ��}�o�v!FTw�\�&�����;#�p���S`�xj�3N�]]$am�&^g��p��XlxVHYEB    2864     8d0�K���8�q#ǲ,�p�-�-���0����kŅ�$��Y��'ێ�~��=r�a�)j
R�k�(����햗7J�-̔]��l�F�sO�v�1�\�����#�u��|��B�?k���P$^ݤ�E�,7��������l�L��x�FNDM�{�d\�K�c�&	;d ��?�O)�c�i��+�V*)p��*��)W$N���)ވ��̪�^q�]d�FK���	�B�y~�bZce�GE���(�A��x�
5У��	� �.���d��U��N޾������(uiD-��7鈡� ��l��w�n�<�N���>d���ܞ�zΪ@�y���s�}p�&��q�w(�KA|��ޒx�V.�TK�h4�1^�O���4�4mA�������E��H�k�o��bY���Mr�R�܄>��,�LgД�M��$7ƌ�-
���S������!g��
�$��}�4��Ψ#/Oj��0����8Yg�8���o��F��R��eG�p'�2��U f��� ��ȏ������GP	㲜�u#^���ؑ�^���Gy��Nn`����-�Ѷdw��ķ�%P{�I��0���?)� Ц����vQJ=�����Iڋ����>�~�H|����� ��o���6�(KT*��ʘ��vA���)�-����<%M�����	ivfb�i��[�ɗ^d�g��w2�;y��v���j���SFǒ��|~��6���N@!ԛ�A�)��i����x(��3w�B��b5��DA�_r;�;߼`ؒ�6rʣ��%�r��RtMJv��0i��P-F������Qm�;�9����2�k���X�l�o}ʱ���#����	�j��?!��|�����)� �3l=��g��ߠ������q`K���ono�N,�>߂ׯ�h�߲zf��T�9���R����@�<9X�q�i�[��<%݉D�*�|�d�e��p�zrrP�n�-���RP���q�ǲ��6�@�1��O�\|:R쑉2ʖ���Z��:���P� ���\�A�b\R<�q�̸�x��	L���@Ѡtǋ}����k��n���E�-`!P���}�1O傭r��,Ng���!�[Yy�~��Ӈ�I�����y���MPغ�΃�lE 2����v,��l�L/�iv-E@EHǙ����)$���v�������K2+�g@279`p�k��'@���,��w�xUN)��Xe���o�u-�H�}U��j��6a�+hkf3;�9���ҮEf(��vX 8��Y4O�/^9@�He�jH����~wJ; ���pbU�$<�P��x�!o۞�>��قIFO�T
{RА戕�S�1�)�+�%l?�Za�0�ݛD�F5WE�aRA��pz	��Т�/�k��O֡��Zog���}���dz��R1�7HDM��� �F
�g��.����W�� �CKvD�͕�->8	PCvk<�i�XJ��S�8'�n+m����&:������g��?��-��J��z@����Ew?���i�:jkM�"��Z~W��<�`���^���\w
Uk��m��+clN:�R�l�s4翃J�z,�U?Q����P밭�+U��iY�&�xO��H��?h��=/n�m]�b\������f�]0��((- �>���8g��"��Bb�#���+BZ>K���xHr��{J4�u�Dv�6�]r��m���M�<Jw�d���ɾ��j�fT[��X^Q�^����>)G�����Y�lj{FڕVIU���F��e�c�+�R�d��"e�~�kj�x�;�� Ҩm�x��+�)=of'�晭�u������$`
^5���}�xR@�)�"c�S�fx���Z05ȁ�W����jF�~"(aU��H&�&�b��a���β=i�q��{���E}J�L$�� ���M�Q[g0p��F���Z`-�� *m�\��ߩ�䲻(���x�>�wP��R��oln0(�Z"������Sk�I�՝ؖ,�L���$J���j�ɖ�@��A���'�I�tT@:e HQR<PY��;�n�YЫ����_�E�P� �*>���6Q��O�絏V��18:��$��0Ep������M-&��:�a@��sY�I斀h�\�h��Le��j���퉶:r+^�y,�n2�9�rЪs0a�4c:G��������'��� SN�^32��Q���	���Ś,�]