XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������;bVp��4fG��O�c*����/h9u�ޤ�]0�O%I�)Q�]�O����j��u��

Eǩq+%�����(=�6�#���KOLQ+T�_�3��
��x�t�4l?Ym��
�m�	�doX]8�w��p`E�S\l��,�>�R2��~J���O�	7|�=���?�!?@o��Qȍp/�|?)r8�Q�n1�&m�l(!U��d�|�6��V2p�'�h��o�ff�3MJ(�5Ʊ��j�c��V�P�MhO_l�p.0����|�h>��,?J�aO��]��y��>
WJ���rY��м�26G�I�*�cCܥ�	��9>����.
�����cԌs9װCTX8�����8�3,X/�N^�sh��h��� �6�NUb��C��:_�J��y��*�T�����s�a@�Z�f���\Qa��#h��;(�I���v.���aS��C����6Ud�G�Tx�j��i��[�x�L��m�[�/�d�MHBJ����ý��a��"�	792`����^�N1�C�PU4�-�k��[�����*�a����c�0�
�ԇJ�9����_t��}�.���/tF�H��\���跢��V�D�3�`�?�&zA��?.G����� �L_#�:����8�
��MT��~'�	��'*�jk�a�����%[� �p����N�Qt����+�4CB%��"0���t��u�Z$���Ŏ`��ξ|�n�ĺ�FN�Ob'�#�Sb��?�:����XlxVHYEB    1578     5a0ig���hAˋ"�E
���e+�qpZ��󓄺��،	���Nd\k�: /���-�XR�n�?/��)43%JUD������[T�xk$��C
T�1��D�G���5<���9�I${p��=bw[�Ǘ[2Q.d]w[����1�=+;�"��*W�5��(i�4�~�Bc߁���|F�%��7���zc��/  �a$���Ŗ�;� R,�:D�͗��=C�Kg�(�o�� @�ğЎ�hM�;���D���z��}���HI3�ٖ+�g�q)�-�	�#o�<:��CY�g�(��N8u���U�v�\i�-�&�2�H��NcZw�#h"H�N54:O���Φ�O���.���6�����~��P�"����~��cbI��,-r�^�ޕ��@'~"�ԗ��������E����eձG.ߤ�,���r$�*xP����NK��[�#���Cm��i�_}pȕa�8�����x�����
�U~z`h}0��'�&$�~p5v�� ���ֽ�ڭ!���@���
,o0|:�"U���6�Ur��	hcX�@4JWP�m��b%�pW�#��q�].�"A�q+�̎���/�ȉ����K��z:�w�v��U�׌�6%��ڼ�����H<sW�L�E��Ӫ!9�M���DH�G�ٜ���*�b�:�. ����,]�����C1��!\��r��&Ư��^�l6\���/Kp+�7M�����\S�@��� \���a���^�ʬ��[td�'�Fu��w�&6o,�/-�7�%�"3�w;]�oCt=�q N��>U�@a��Ǝ�0)$�B���7W9�@���ˈ�mU�(�I&����S�ׯ^�uw��~OS9�� &��,�af~�`�R/�KuJ��<�Yio\(��B���+��_���	�Z�!�F����`Ѿ7�{��Q��M���cD�[�ʌG�_�񺇌��2���'
��ЈhO7Z��̦Csp|�+�Ye�v��B��G⊱����ل5+.����;3F:�1���z�n_~'�
$��a�`�3A�X�Why��B�N�\8��7!D���r%���c�S.5�)���=y_��H��	d�������_QA{���d����c��V��Ͻ���1ϭ��~w�(]���OY��ěVOm���6rܗCV ��^Ph$�k�N�Ϧ�R��\Ul��G"�d�@�`��)Ū4�s���C!��K�ǹ��6[WY^#�ֺ~0X�G��4|�DrZL��{!���y!&���C���O�T��w��%��<����o�瞔��Y���wo��I��D6
:�Vq@[`���ٷ�o�0�5���
�*0Ru�aq�g
�Sd7/�r��-�o�r�w#�J�����$�礸zK,��È