XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���{����{[���8N����TQ��P]�KY�`d���7��}�l-����?tz|�Ȟc�I]���?���t�.^��N���p�Jec#?.�c�80��}�������� �W�<Y���m���7<��{^$��I��e���U,ud��V�c7	rJ�Xp���?�� �t��jO�@eT�Y��*&+L$$�)���4�`�e�z��!ZDb)���8ԁKt`k��b@���K�g���ͩ����Qn(~(:{�� flX���sf�0?�_��P8ŋ��Vno�h$��Y�n��	V��=3>�؞��W���w���9�P
~]�2(�z���Jӥ��t\�ڊAʪ������DL�_��j86���c� hIc��J�m�u䲙@� kM���u#C�C+[.e��	�Z�a7���x{!=hX��"!��v�Z���~�u�R+O6qz��[��11�QBF��\�h�k��ɣ�G�ُ���l�.�M5��''R%e#�5;|��\��DQM4jdL��B�٫�-g}�ظϥ
��eÇס㬽�b�SH%��#v#�]	i�a�r�&/U�J�*�_4�x�q�
�N�R��*���
l���u��p��!�=Ö���SfT�����b���_��L�0P�e�<�E���o�"<�<�6�,�gH<���9^���>0�'�]�dBi@ȹp|�_�.��w�P����ϧ-Lg���Ib�]�s��K{�c�����)���?:1W��@X49w�XlxVHYEB    312b     7b0T�Pч�i@Wt�^���4 ��g�C|�ǧye�'_�)����6�ӠLJ�e���t����g��j�VwP^���'rՍ���p�!���oз����Թ�r��/��Q�߲-�x^�s�o�X��!�M�t6=�k����:���oa�@±�FK;C��9�ga��7j�����Z��$PdA��X��f|7-�e�s��
����"��ad;u̓w�T�M��i���N^�w/���u�m+cl��\���F#���s}��D)BͤZ� jw-�x�X�9Y�,ͮQ��q���ǹi�`�i��k��w�DD[p��W;b÷��6�N�_B��������h�*\o�D���4$a��ax�m��c<+�fS�G���B��X1��Ps�x�D�b菾�h�x��� -�8ѿ�(r�UJ0���IiL��iϦN��8
<F΂Sȍ)����X���4@I`nG=u��Ϯx.��A-�`X�VNjiy��H��73��A-�<S�h��tS�ž�du1����#���$���=nc$yR���2�ܳ�ɨt�)H9�؊8������1E����|�*�/v5�A����ds�{����(��"��q�?�A
�_H��
��z��=�X�}�kt;&@ ;X�)OQӪ."������Q�C6��,��6��&�����y'm���� �h��g��{��)~:�N�[z�+'6�H������_���w �/ԁ�/֩<+yz��^Y�crP��d���B����:��קl:FU�Ii��'�(����8����%�#�NƫC�o��}�C�t)7��l�z��E:%Fw��.�~�C#qNz��`㹆�Q�k��芙�:ጶY{�#�)h����m���y�##`PQL�ƴ�B�27�?��B&��n�%� ���ǿd��sU�����1��@�(Ш�K����3���55��Fe�A�f�u�m�J���d��"��5��%@������%�Ky�?5�jN-�k�5�����}
>����[�(�;�J�y�J��)4ʱ�����MlƬ�!�3h��k�Q�;� �+f�S�1>S��}m��ɣ�E�TU
�q�iw�ث��X�!x�u�Ͼ&:��p=;� ����g�����,x���`-mM�w��>|���F��*�a|�1�^ݲ!��T�.��	$ɏ�p�65��T����#�|�nN:�1	�p8�ko5���Ȩ�Whw��,_�����o���N�Bn��ޠpa���,ꉡ^��9$�3v!~�|��!Y�.!QH��0ᓌB��^�>?J��"��jS�;��|�ܷ>@YUZzM;�FS^��m�i_��� ���3a��ġa�/���\���'_��Z���!;Ʒ-}KJ�@��V��"�\
������6T6�bH��#+��-M��B��r4�>o��_{:���3Ρikb�a⠫�+ �d� +�C_w���<��&������*�_O�؋l(�Y�V��Hzɥq����-��>�"j�
g/�+[��vH��ߝ(�Gx<���VY ��G~Eq���0	g��5�nY��,#_ɻ�u�k�|��`T,��e+�w2N����ڂ�Oa�1�??���k�x�	�A�������5�:�FЮjF��ȕ��4q� ^�0"$��.��,B���@�ݗ}�=F�.��0���"�8�
ݕ�ˡ�T�{*�Z��ͮׄF�*��0�w�}֚��I�*��O��֧M>�śK����n�Ȕ��?�*��t2��aZA.e+B�����g����6+��֖��<�i��a����������Yu۔����2�v�9][M�6L����J:��ֆ PX�wTc����MQ31�5��"Ϭ��o�r�) �yL|;�?E�\(� �G��i>K*�u�R��d�5)�|=�<� 4�ԓ��y�Z����j���L���9�S�/ͣ��L���]t���