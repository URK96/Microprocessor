XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����"�����A�	A
C���Ռ�o�ZI:v�h���W��b>���rBeB�B���o@2�DQ���0�ӭw����tGZʎA/�o5��q���@C~/������,���S�?�#3� p�K�z�X][׫�@�cz=��p]܌�s�$C�*t�م�>W-�45ّF ��h�C�J�2m�^�V�5m�EGX_Q���N��/=�e�I�5���B������;b�*�ʭ������(R44�\E��a��O!����~���)�"��s`K"�nJ��t����Ы
�2x[�- k餙�T�L)-�4j1>�-�}��B!�A$9C��-E
ٻp�OD�I��W�:e>��S�OF��-����_�f{�1���ȀL�Ҩ����h��,�VT��v��j&ݧ7g�
4��f�X�2��o�M�b��q)7, g2 �����y�;�Oۺ~���o��w����>�l����GD{鲮�R�� ���k��V|�?H�pjHiEd3� ���"�jv�fp٩i��>=���@�s����5v�q�v����U�9�n����Z���g����z���J�G���/�%2�� ��E�i)��ܧE�1?Y2h|��ֲ�r�{I�9�,��AԈC �ߎ�خ�,*ߪ�?P��LY�D�Lu�
('E��w^��o���랮����
Hr�e�Xn��p�/k��;������N�c�w�U�L��y�+:_�����a�BH&�XlxVHYEB    1001     490fm7����ɐ@���/X0D���n��������H�wi�@�B��7�	V�%/�5�)���S�hAUM��+�s�Q-9,���c'j^іØ��-R����`/>���9��'�'Oa�HϽ�P��a�~AZR%#���4��M;e5��c�Yw�|���k�����$�T''�cS�w.2d�M��Q�cx��>��C���tm��`T�~�8X�#��/�hl�х1�ZT@'.��i:6~u�ԧϸ���0zGR��IJU���f��A�.g���_VO8�?�x�[N� .`���<]�%���S mv���u��W����4�π�́T��Q���aZ�sA,��X�������|�. �4��絖r�K�?(Y�&;�4a���|v�.�!b-Y��a������[	�8V�@���(#�`L~��pS�5o�EȩW�����f��+]ŧ���T���a�bLe"ʕG I6r0�D3�|���`�����'�#�äaab)��-�❵<�>�ty���ݩ�� ��oΔrBS���d#�eZ�
O.Ѻi+U<W�՗Mn�f<
�SL��4O"��z6�����@V�0IyM���C:4����>@ّ|�{bG�[{ ��&���r$5Ӛ�5���W�CG)�Y}7�"ŜʑM�F�g1O�����k��sT�� !D�>�.��y�,��]�6��4q߅^���z�xvx���=��B�.s��7N%d��|�n�u�
��~��u����G�ِ�IήY�����_��iM��G]n��>Z����n��c'|,�P��Gnb�Vy��2��0��q���'ˁQ�鹔{"��
��:9f��V�~R�}9��^!�U�ъ*7��Gw9��[��x;c{R,�T:�?D�w�a��wt�t���-�$Ei��p_k��WiA=�����{e�}��.�K���9���u�F��i'�m��:-/����zpu{���k�l�|��-w5�Q���!~�X�W�`�`�Btt)	��C�=� ��I�H���Vܲ������c�9��s5ĺ����f��x�p�}����t��UM<B�Ě:�<�f������抴k{%}���i*���yV-�AL<@�̂��M0��Ҳ��4��"���