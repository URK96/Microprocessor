XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����^\#ܷ]�Lo�3q���?D��ÿ�xD�Uj��R��2�QDh_[ڪ~�����0�e���_8���c�3��k�<�p`�Jj��Ҡ�4y~o�6�u�/��jv�^�� μɨ��	��9�5	a�`���
8CjeE��,]]]����d�p��#����?�����]�j�/��� ���pG��*	�Ɛ�wZ��^�\�)X��� �A����R�G�&�0�F{��:k6��:�5Iɸ�y ��9VF�w�ź~�t�Z��#{�K���Ӵ��Wrk�C�0�vrn�8�g�5W�W6��R@ś'��{�a%mMgdY
�Q:�o.�$W��
�y��P?���:%�h��Yv���0�F��$� ��?��äD@߀Le���ͰA��5��Q�g�`����t��0����s�W�K�#��֒H��������+
�Yv���-�1�?�( �x���8۫Eh��+�&��[2����v�	����lٚ�"ի��1gj�+Q�P�6�eQ��cD]D[6Ӝ[��a�"�?aǈ�s���極x%���<�R�h	WWI##���Ptp�l.�`� �ti��ڸd���u]<KF�X~���^�ZM��5nT�����a��� K,51��<�p�.��[�n�yrLS�2(\�ƒ��A��8�/��M�a��0Jb��c����̏�,�� �}}�ICP]����\w 5
%4-�j�,�Lĳ+�P�2���ZTqb�'8>D,"Jn�P�(XlxVHYEB    152d     580	Nv�:?~�#:�_�`�峷���чck��#s�er���Ԭ�h�y�������G�A�|Z��X77�l�܉%�fK����9.�(�p_�${g�΋9!�[`_��e������By���E�v�qY��i��PW�O�1Q;)4/؇u��U����h��~�%�i3L>��k�hX8c#�"�q؂�aq;⾝R';��$�g���<���,�����\�$[�[���wd�볺 �+�$qo��:>�a�P��o_`q�Z�wE���.� ����HΗ����]�z8v�t}	��\�9�B���r�)�u=Fu�k��O(6��s���wm,qT�DM�0R���[�4oC�1貧��^���k�U�&F/]�p���SC�і��� � 獣9�2�;�-��wVƟ����0>oZ��ߵ8^�,�R;O�oKEM v5`[���;��Ib$|CaS��������5]\���9��=W�XM�2���^9�"U�L���f��uK��~�BqޭQJh���Z��8�i�R��;�_����LӸ��LF��1#�G����Ɓ����T�g���[�T��^���55�N�05�3�9�Uq�LjNb�y�Z�ˌ�H��v ��X:@> �nob|V��I��ce�}�~�dG�!�4�e���|��NoŹv�]��jEH��M�z������3k�{����K�����������|�%�,�K��/l!��V,Oz��SHMG���[�_��f̟�F�rc�tZs��lB���m��&O�R��u�x̠ �M��Ag�wu��y���Ts<8�u�oG��&<z�ՖS�T�#Y�Y��D
\+u%'������i�E��p���O�u]��?�S�?�c��L�ל]��=���uGe���Q�#O��6�������o'3�aI�ɵ����V�S�j�)1�'���[,��������)�q�U.:��X�����Y����Z8�<]7��`0��g���g�w�R�U3o\�=O|�D��l5�w8��̠�Z5��f(q�w�ٙkH70�Mn��A��k(ݼ�*k�Ar�B�M�g��\T]�>�v��П��f~<�y�=��{bSn�h�B�
ϱ�W��>�@��Z�Km���!���5 x}�3?������J�e"yAH��x�VWO�����y��P9�ۅд�dP&+��:��QC��Nw����/k�*��K�J��h+��̣$&s�)�`�Fk��C[��3��s��1�s�ь�Ņ�ak���B�vܫ��j�7�`b5�inҗ5�TL �$��/2t|��n��eܿW�S��o��la��6��Uf@����?���L�ꐢ�X�]�~6�Cy�l�xjv
x's/<|�6�>�܍ݑ