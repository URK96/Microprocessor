XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���KƮ�" g�	«���݉�<�<�|�c�?"���R5����zy����t
�B{��ҹ����mJňg�oA�̓p�@'Wk DC�_�::#Y� ��O*�/�P���Y��'o�G�x�Z�gL��x���ш!��Sjase�� �x�����?f���!��$N�jK���y�Vs���_O����C;2�^抹��
�����mU+h\�|�Ù����m`x_���-��d�%��9 �����\��7�WV8�ev��93�T#+����L��_�{Z�-g`��Z��A 
�-t�կO�J`�i����dd�H���eB�i�/��vr��v���L��Z���@P�S�_����-��yl�<��P^�N+����F���fJNs�>�Z�Q��4PTe����ID7����%���
?Z��Oi�F��
k_���A̱�\��
�'�%J�hI�	�k�(Y��?��qE^��W>�B��_��\}� ���I��C��@��6��p:&�[����sa�Յ����9���%%�I��0�ލ��V]-�s��P� �kU�8c�����V}�]���S���l�"۬/�f��ڪ�+�(���c�&%�c:Q��m�f���$&Ƙ]z+��2k����ւf�g��Ag���+V���[�MT�/������R�o��2�Ҩ����R�ϖ �=N+�9:��o��:R�����Z���;9�)����>���!XlxVHYEB    6faf     c30� �h'G�'^��{��ts�.i�S���3��r�4b+���X���m��@��0ڰD%Q�����[<�?0^�Hꝋ��yCВ��F����ަ˺>I�W�IwBQ��͛Uc�>&U�kz�Ks����{���.�M�|�-��C�+G�&eI��6��#ŽFw��l��sկ=,ʞ=�]�ʠ?r�Jz`�Q�璉�y%dB��/VPWE�(8�}]i/�\��6������aR����ET��g@���$���ù�\]�s;O��SǺ> f7V��?��Ft�:�oK����{��ުNh�es.���Y�ݵ:�5���ю}Z&J ��n�9�s�u;�{�yg�,��M>&}�&I�袴��h���S���m�5DO�O@Vg����L�u�2��]�?�Y�孢�� ���n��ky8�5��٢�����aZdP��@�#��a��7����Ø����xR���~��o�ǐ�6<Nm#/�zkyL@|%l'��-N!���� ������� =@� /�Y&zL�V�W{7�3m<��$*9h�����BP����o(�8����U_ir"�^I�`���y�����\e�G���b�07��Hq�s+�ӗV%�o"�_r��S9Pn:���Ú�=6uN1����HUyќ:� ���+j�1ʛ�T��QL��~5�s͔�l��[Z�;��4
?�C�|'[�cgb ��	؉�t#��1d|���x`��n�$��f@!*�7�̩4�ZX�ZK��q���CF�%.��k�a������p�.�%�:��75"���t�Q�HF���M_g��p@pܲU��&�&��_P>Dޣ�C'���O�(�S���5��.��I�SvO7�`H��=��s?KA婻��8b����C�$����Ԇ��Mŧ���oS�:����KM堮�i��Bx���
\���;]qs6����$�q���%N�wԺ�RF!�,�����s���n��jL|��%Cҗ!��փ�Uҩ��f�c�<��=D��t�G!	>\�D�)?��pDm���eE������&?Re^Gޛz��P��޽8*�<�9Í!��C�(�y��$�����woz4�wVp���O`X���nK�-��ܗ�:�o�w�y��C?P�1ᮬ%#V/:y\�	��WVG͊C�i4"m�4�A�3K(4j
��x�9_�,��+��[P�1��B�V���z�����o���9�0��"A*ȓ4{A��&b��K�V��lȼ$b���j��e�G�� x�z�ԢK��˚�����d#��$SI��/ꉍ������ ��RK�䘁�������5O��7�x7p}y�,�l�nҡHio*�GB��]��u��Q��^���vf� ni���������T)nzOl��z�ۿ�M	�F7�5�q��D8(��� zo����t0�/v�ݚ������exK�˱�T���Lb+D�}�8Z�˳�ຩQ���r�\���.�a�7�@?������7���.�>m;z�c*��k��nyJMII��}U'��r�,�R
"����ߒ�h�	��x�!A���%�Fs�2�͡n�{�0��[97h��v=��%F�6,��yG�Eh�e���Z$p����aL)`=+WR�Y���)�9n�M���wA]��ڦ�e���ZL��ZZ��\�=�`�?w��h����!e�v?�"��1��ix|幎����Bmo��@���g�^�1�ٳg|�.����u!���_y��m�`� G0��*�Um�dnZ�V��� ڙ�	J܌��:������di$�up�¸��P#��[D��������b���	�+�zhbH+��jF���8޳����Q[��������űS���@�pl��(D�/\w�a~�"�;��]&�f?�C0��{�2��ԧg�b��by��Y0��e��~�'`��>s6��1�|��B�/�O�6���w?G,���w-uk^��W�$+2���i�w���h1�����v�'��K��$�5$���>���0�X�L_�(&"w��¿2����cm��$:p����7����5�0�۪Ώ7�d�����h�µ�9�1�@�����
�Bf'T�*���Rٟv�X� ��J%�-h���C����rq�����^�W�Hoc�����p)����|�l��DO6OIٸx�5�>|��~���y1��x�`��j����8AwZ�X=w:���qǺ��c�~��;X�:��Ƶ�$�5�4��}�� ���?8	0 ����q��?��J����c�vX��x�Q��Oq�쁄���{Px���%E�&��������ZNb�v��o !���^��󋄕�D����$KHU�>?�No�Ō������
�n�G��c"Y&�D��<���5�������gqYtzox�a�x �4�M'�D�Y1lk ��q��Qں+z��M���P��.�!u�.Q���F��PՊދ����|��x����W$��O�3�#!�b3��%\NH�t�5��B�r_U��]vWF��X���l�/D�ե��6�!H0�]T��=��礵��0\d:�ǻu���Q�P�=���@i�}�])U3�%��^J=6����J�꺚��m8�cD۳�D�&")76��ܐ�u�\�3u)g�l�ғ��&S_��Rۧ����hq93��Ѥ���z��'�z L&,#[�~�7�t�v��:Thp�Z��Сڔ�{��a_K6�����lU���=�z�!�z%�{�:ۭr��l�AT�ҧ����o����;�'��w�l�K�bx��F�~�/���;��VD�#�k�@o���M'�ik�������?i����'���9���Ŀ�T��?�Dm���1�e�`ZNq[�EX��צ�%�}hp�S��� �4�Ղ�p���W��D�ք[��<�v�z���3�R胱��O� Zg*�|{�-��ȶ� �������̹������ya&�⏢L�����f�X���:��OۧEC�d�ᔠ�g�Q��A)6SB����哝��o