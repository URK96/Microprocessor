XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������˵�I���P/6�e_2�|Cu�K�g��I���C�	[��|�P��+����Xk� bX��5���$��ߝ�Y�?'��~;� d��eJ�k3���+G���y?bX��W�vD����A@ȕ��-�����Ba_�:Kn�n��\l�{HY�7�Q,�-�5��q�H\�j��r	R��U-BѦ 1���d�u�V,�ߧ����X�r!���=���M��w�r��L�l�,�H�O&�ft�����U��h��H�t�
ne�����A�	�&'����~!��V�קF;.0OFbD�����t�� 7���9s?^ ��Eח3no�y�WgS-q�d! hTܣ�^O<?�]Qhz�}u�}����_7k�+�=���Q.��cxa��g��wM�>[�Q���C!`W&r���ki���|�.�-��F�5���ӝt$�,2����i6�(���L�C7��(JJ�c��ΰS��9�Aq���a���8��%g��D����}hoC�;�`u)��' ���WO*/�@�����7�L��j�
�^�6e������9m&�D��)}�pM����1�i��諢�I{��{���_@��T�E #��u����3�������/�M6�P�KcgԌtϋ͜�F�x*����T:�T�VHG��:lđo�t�4�Y�w�Ǎ�u���_ >B<ۺ�8q_,3#Q>�"�������@�I���0�F���a��H��"okvk��9kT賺�6�9��[�8w\F�XlxVHYEB    690c     b10��oWC�	� �W�av#"��9Il3�G"x��t�bs��H��Ӽ]�f��nϽ���Ee��}k>�Q�Y��E#��Rlg��l���X�M����@�
�]��,�K�j:m܂�\� ]ĲD�_���Ĝ��e;jm�:�s^A�Ԙ��%�KɯN�����j"+��E@;���Z�y��6N[�X<��Mk>��m+�K[����'�W^ս����!��O�%�P���TJ��vF����mCEϫ�����!9>���5��Pq��svl�đ�^�\,v�Ԯ� 2�cC��.]�k�S��O�$%�)��2<�+��u�Fύ'�Vk��z�H��@䖃���z�2�Ⳉ�~�$���e����(����9��(���$�--���$JF�5��	�4�b�x�Z�O�C�8���<�F5�;} @�纞l̙[��]BT��:����T?fc��J��ID��h섨+�4<+?�<,�P{���D�z�o�.�5[������뙼���lPnF��l�t�Ȧ���Y���XJ��G��V��k4@	�IPn�D�i~��}��y�;OW�X�A����.8�BЃ����9�mxv���lC@�a1�e}���)�3��˅<��2�=�}Ӽ�2�u�kY~��#/rw6��K� c+������}���� �rin��2��r.�����;����`Q?��{���6 �X��{l�ew������lno0	����(����PX�C/����Z��*ł��@�9@�0�[9��e��f�A�%G]��6��¡�Y��|/-jH���s�����K��F������th�a�� Y2P�:;�M��K� ~��)h�?���'�$J_Ò���$J�+C����.� �R2<������elI]�q7e�-�E,�K���G�V���\����(��s��Ú�gi��42˖ó�k��W����8!wX�:�@_��#,zd#F"�B�S�m7h5�Z�<��*��;KTo�@H��\���v��ז�#�v#N~��ȶ#�@;�÷R	�����!Z;e�*3�ȩ(+��?�A��[3�o'N��%	��*�0B��N��]�M���A������C�9|�Ws�F4/Iَ&�j����9<��a;??j�1~4�(@�ܮ�KDW�d{ӧU7�,�$���N�᷄-G,%�m<�dk\��G<�+d��_������G'�N츋��O�������m�Ǿ�����xǱjRT��<�ģ�އ����zla��Ƨ^��0T.��P���
6��;��uAu^C�m�G����۶�oq��8�2�� ��&.c\��̫\�4��"9����Zt5�E���I��j��al�sp�އ"G;~#Nv
��G��x;~��g�0�W]����u(ߎ�T��ƪL�n����y�VYDt�E��3�#0Ap�y��-���n��ƅ_}F?�&�͢0���� ~��jB��rn�2�+�+|Щ`��3:%�]���G[S�m�T�g[3��{��n������'|�g@�^�5��\��ݲj�лu�kB�a��/���d�f.JY8��%���K䕿L괒��X�쨗�s}��e�Yc֌6�1��P!Va�׆�O��'h��s��7��aLԂ�_���zmn��'o�]�"�W8��{(��<��_� o�S�x}�-�n�\8嗝50Wպ�'���HB���{��u�"�2vv�oP�zB���>�Y=?��M9_Q���8��`�H��է��C1�"��d�AjX�jj1�$�� �Z���a?�S�5[f_F�	�7��%Hɮ5Ƌ-Q��H#�� ���W#�y"��uL9�/
I0ǭV~�*K���&�e���|?H�1J��5X�P0������W8�	�sڴ���Lg�+%�N1����>WkǺ��RTZ�G���(��}�褬�Ú5O4^ܶ�8<tY�LE�*��@I�� (:iUqAW�n4֡����N�3V\��p�Hh}܂@�D.n'����j���0l��	PD�-?�� :�مoy�頜���_2��'0�|n�K�r,췽��������p)��r�gM��$�e�r��?�8x�K�S
�f��V�#������pE<��g�%Eݚ�9�'m�n��ʹ�el9f����8%K~��熌1�ۏq�Cf��-�r��rP�NT��Y�G��<���_x2��<l_�Y:׏�}�*2t�Uf�2Vn�-O��;eㅋR��"N�1�"ܢ}�N\�=��7�f����w*(4W��	�x��)&B9��r����c޲)O�S"S�}}��Lq�;��-��
���Qy���
k�͏����>��] �5���{���Ȅ�UL�3�J$2�X�e��%��IaZ�<�t��`c	��`F��}{�͖���jQ�B�Exc=Fh�@Y�p����I����:�gU5hŨ���� �;����U=����vw��N�Khbeߢd�Ep��Z�"�"ֵ��QX#�/�ϧ~D�U��H�b�[U�m=H�Q4y^�/q1hQ�Q��H�Q^Jj"J����\/�e�37�'EK.3 S׊�Ӵخ���:!��~��o���rw������z'�qs0.��Y�����O];R�L����[=rt!eJX�NW{�M��W�'�9�� M��VJR��.�׸��ue 6���ֶ��Xݓ1tt�lw��4�ǧ��Jզ��R��.Q� 
?Q�(�`=L�j�	��PGoCT�