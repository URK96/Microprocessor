XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9�%���I��������)�Aw�2�:Xͪ�!'6$�I���!/����H)�լ18��b<Q�y��2b ٩�I|&v&\�u�ؾ
zb��� ��Nyr�]\-��+��k�I����E]�vVoE��ݘ�r^~�(�CJ���z]�EDp��uo�_�|�D"��g����p{�涾�/9�{��"��w���h��������4V���}U~@HwL0�̡�?�&��z���u+��<F�#\�}��R|&+����pL;P�z-��P���&	�LslN��z{����?��,�r�F�����M��]�|�x��E����HS@�FTX�,E��E
ь�Gv�(��}���W�/G�uXՀ�_ne.���汁� �`��g��;�',!F*��:�%v:��tk���H�_4�-�!��O<<���$R�nN���H������8(�q1�Vq�_>�P9��O����?�\��E1�R	��b��<ֻ�ڜ%f�d�Vw��}A��?j>�|���m�� ��Po�������d�ԖW�d�vIw��?�(P�&ߏZ<�5�W�e��qw��Y������T��b��h2G_��E���%2��Ś��{�G�w����Z�k�7��-���V�[d��][&vN�5M~��Di�.(���Tۿj1�y��A4�8���3�	�w� �3)��n��`
�B@��Ⳁ�6�BAb��yie�[��)��qs�>�����GxW9XlxVHYEB     9cb     230-�+,3	ŭ1��Yu���z��,�ANU�9{��'�jG���G�#��� �蓙&����G{�o�;wn�K#c�p�Y���;��C���C(X�-k��MvP/)�N6��ʹ�A��ᠩT���	 ���nj_� O���ce7-���E��0��G|��h�]����ŃN��	¬An�g�{�ź,���h�'�n�P%p��:��U���:�ҍKޠLڭ��"-�Y$�`��I�q��C"��G��r��2͕^�8g(�����/i3;���	�c�X@� �\�G��r���T���>��ۇ��۷ ^�}ūh�X�?���aX���@u�h�ی7��uҰ����$~ī(�֫�^�ǋ�lv?��ɸ��y.�"T{�/��ow���@vK��A�0{R��I�WH��X�{_@�:`
 ���;�Uk���F���l-�3}����Lj��|L�pY�y�w��@�� o�,'��^��`K�6u�����2J�Oc|P/���}�@Q�Os����p�
�{`���X���G 
�u4���