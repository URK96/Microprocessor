XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I��F	a���s�Z���q���"z�{N��Pt_%�E��T�h��\j�w��o�c	�]�Bdt*�߈&��n��TAc.���NI%C��Q:�/q=斡g����t�?H���܌��w�� �͟>����;:72���w�ng�}bݲ�]Ň���`�_\�&I�ԕ%sd����LɁ��绽�ð@�+C�;o{D���s�ѧmB���*��08��{h�.������=�sQ`��R��˰#S�`��ou�$��/$r��)#6�K-u�4{:f�,�l�n�l���,�* �\���)c�0��V*8"�Ӡ TM(�n_�zQ���.�LQ�MqHg&�|�_!L׹[��E{ݩ��c�q~H:��
u�B�0��'�d�"=h�K<&�`���+h.Q������2'�w�:�+AU�á�h�F�`_����G߱,驧����3�\��������i

˔$�9w,
b�eց�.�yIZֹ��f�� �� �bY�z��E�{�a�q�F��WߟL\�+�[��1�Y�|�z����]�2�ҿ���>M��v��"L���a�$�`���5ތ$P�Zڌ˒��������L-�e5.)l�Z<l���v���B�^�� n٪���v�g/<��d)���U�c�B�W�/��S�M�g}4��A���r+�^��C%Fe������H�0�p�� �翎ǘ<�����Ş��p��EdK�J�)����K�1���L�#��vL��P�XlxVHYEB    fa00    1a50F�,�t���~�?��;<=a�-;=�o��L�|�t�U���g�_A�Vk�����K�JB�b��o���؜K^N(A�"����.�:�WRĈ�Q!�셒�Cw*@���@:QDzQ����WW-�X�}r5�^2�/B�)}����#���C7%���-�*��߅"<�O��No+[�#&#��[.'TR��v!ï7@-hj���Ty�Q��3�XG�����vC������'�q�J��6Ψ�*��7=�R�����	(��֤�	8O� m�ڝU���Z�0N���WNɂ+���y�)���j�F������t_{	}ɠ�:L-n��^�����M�B�NW�GҠ�~j��0���M��y�|��	w��S�"���$PwW!d�2L`�n�2� �{�6h��eh?��U8#��r�ޤ�b�_���@b�ِ���@�E#�=�|Q��ۏv�f����"i��Uz^�a����Nz��a�hnp�e�ơ�$5E�ߜ�A+��;�VM<���>��F�n�t]Jo��7�Q��"�Gbđ�C���T����ؿ����8,�O��dqg�"f�J����Ɋ<�}�˃�׍k�!�;:"����x�7�Q���`���ۦ���*
�a8B?�U9[�\_�7Wۚ�|D4<�L�]��ǈY�n����1<_n��z��4a8_���k�h�Yt<���/��P�Į|F�&����7y?�)���9������E�,��C���K2���h�����X��yM�<J�f�0�
gs�c�l.܂o6��0�RV���<ר���1M/���~��X���~Q-�C�k96->
S��vI(1�c�E�Q4��:�~�L�m��&�X�F��'�4�5Yu����
}�1'9�H	c�$�7Y��X�~?Y,��~\t���MK�W~但���`�9�u����z���asRZJ$�����e��Oڶ[��(S��Pu�������]j2��EO��D�JO|��E�j���[J,"�f�����3H�yS��!B:44d ���_�H��1վ|c�ˡ�º�J4w�M�_��yku��9f �i�:AX���OYv�%��Rzvؿm`EXba&Tشy�jS�lNL�d1����{��_G	�ȵ�r��z�\+��ֺ'�R
vQT�AM���Υn��)��j��v-k�0�)������(�	���/EȤo��-���IH��<�>yR�Z72�(G���p�e%�l�2��;�xJ���͞��'j�
5�� ��)�vP0Q��u�<W�j����A��� ��0�]	�~؆���JHwe��噖g.Aҁ����"�����ʜ�T(*��IӤ�#���,\�E6�{E[�nǳ�F�N�!˖�$��ޚ�Ӛ�y�ޣ�H��;O[�y{�70����ӟ�ޠL)��m�n�E���� ':��a�'MC�ኖR���߀�G�/nf
"?z�uM��V��4!2ݽ��!m�Q��~Z�i��P01�֨~�Y~�CQ�\�a��2�cш��H>w�볧�쳣�^��6�99rӹ>M��gE>%+�[\�����Ҁ��au�Z6��r�m�OKa��{ ��E�.O_���j��m������MPe&��n�	P=0k;����vqQ��1>g2�8n'� 9��@��c ����e�%ΞrC�ox`d���ZG}���l�*������j�D��&�J����ߓ��HV��F�9������b�3r�D�s.���2�{'�t��T_����L$\�5l��b�v�F(����U >�ڽ�}��<�>tB	��KB�����0��P\R����NLi��|6���a@Y.�S��"�X��ZxE*N����<3�P���pN���߹�c�������"5Q�۠�ك�6F�M�_���:��Ҿ��	#���?A��8n���☘N����f��87�ss���>V�ڿj/�JC껠�e��������%��቙2^��á�{_��� K���$B$�PԶ�՚-�S�j10pu0�B�Qe��k<SO0�ݨы*��T;7��l����~�\]�KA�T�'�-�;Ӏ{1[�g���w�`㿻?��u�H;���'�-#��6r�ﳄ*J�=6��m��c	$mRޑ#�Es[�<�n|�wnu�L� ��� %%Ag}�g�Rx�&x#|��� ?�}����I�V���cJ�M�H��ϩ�k����I����XY�)\Q�#?�?�[���xO�Ͻ����gOZ���<�)�!I叝P������2(�p5�c��7�L���;��*�����%��*>$B�e`y�ޭ���E?�i��:g��	��"�0��D!��=(���/ҽɠ�xaի��	��|������PC�ۂ�q�c-�Bx��Y���\m�5[���X�DA ��������x'
��4�t�@���4�.5�|"M��k
Z�^ASb�%=��C�%x@��[(>�Ӟw�pN�pc'����j���)�9�j+6�1�1z�~5-�T�s��12��j�݁��T�kg�d�͋6�/uTs�{y����_FI���\\�0ϵ���xrx7l�ZSWW��_9��e�o��!�bma���S�j�^�� �t+�L���4;��;��wPv�G��D/�.��$(k������t�A%W'�y�{��ªEv%�}�w�	Z��24����@<m�k�j?>���	��Zn��CzJ<���屉O��(E��'c�1�D@��5��ڎa��]n{ⷘ8[�첖�����I�;��2�Gȗ]U�܄��Z��LF\X5��"�S�(�Ɓ�̼/�����4�:.�sZ[��%�L����j<���M4˭���}8Z����Ne���	�9X���J�g���l-�IfT?'9��F��b&R���#\,0ZN�U��&��)���\�G+��\��!Ca���?�V0h��6�����v<��(�kΙD��R����S���~?��4Q�A���HC����>�uH(���@r<��)BwC�[��]I;�u�Z�Pv���V���� �s�aU��=F���ts��8����h&���U	�jD���x�7o�b$�P�h"Wl�݀�lQp|hW��r�M{TcL��n�a��a���*����+��s�'�j��[�Q�rW�J����l���`QK�x~]�A���B���#�I�L�Z���ݔ�C�PŘ��.Y>|,D_>VY�j��%fh~�bdb���P��lN��n.��!����U����"�S8m��m��yN�ڋV��v��oQ¨��.�-��٥�ʡ��ݯ8@�*�P��5�K.���&��%w�0�~;�f�@�TR8
��z��Ǆ�g�@�e��y�@ܹ]�<��}f�(���9�R'�����=a��h̄{��<sPشx"f,9Vü��Ǐ�˱He[�p�j%*�`ҿ�C����(�ҽ�"�����ыݛ+{��7�I����H#�\0�?���F��1�|��N#L�����Z.@nHɘ�A�vgަ$��ڈ�+�RT��8/]��k,8K;	����(M���,��AsÖ}��X��;u�Lu�:�H!V�	��f!W2plЕxF����~��S�ꈆ�*��G�4r�]�FC̄��*F�0������@O�R�i�(w��!/t0x���'��vhB�B�a��c>�����a)!5;����A!�Z�Y��I��D�m���oE�Ӗ�������#{nL�wJ���:gw�pn=��=Ѕ�bBkÒ4�߮B&Nu�g��e��V�������I�)�jm�������y��.����n�o�hQ;��-V���VKq��� a�O���C,�)���,a>&e���.0[�ė2��޳.�>�q
��%��io�8Nqhoavv��x�i��m���VNV�}&?,�ӰNe�7y#Z�7�C�p��T#��{�U^α�K�*��A�)�y�#�8#�\�� ���L���Cw��I��v�l�z�q��#oUy��� w���F��L�s���́��_����&�\k��u��8���ٹC�V�S�Q`��c�Z�K{N^3I{���B��xLЪ~x�v��R�SBFwA�P���E����7�����k4ŀѹ!L��4z��.�v�I�o����e8Qm����?�ă�v��dQ����D�re��5-h���Q�##. ���0W7G�o�%K�&��r[.,�*G�`s%�ij% �r&,�;����x��{4$+
\}�5����%��+�g=�]B$�ޙ���(�	��c��b��^�N|--w)l�~:����I��R�f��2�.u�Ju�Ă��O���g�m�7(҃����Tf����	jV\���2��@��L���nN�D�>��)6�p��䕀�-Aϟ/�h���Ã���?��	Ҁ�����uB�`�ڴ��-ߤArG*�>�}��Aw�X5O��\,�_�<%�r<�O0L��7�w8m>�)����Ŧ�`�dYQ-�RBˀEo"�����vUa߯u�H"�CW1��Ax(���0(��-���E>w������{3�P��;������JI!}�ӓ���"1Gܰf���׿+X;"bB��E�w�:���W�px�2�[gِ\CD^�K�sB5�q �>�6�\N8�|���ڝ<G���e}7�a9=������`<����"R��ƿ�=�̫QA�,��m��_I�	��ڳ��.�� ��,��k`P�����}y炚���b�?���EU�YcI�>�˞�����:RyT���H^1�ç�����8�(sԊ9�f����#`D�k��f���Z���w�a�b���˝�`1�4���}9���`��|�.L@`�t�L*Vܠ��\�Uv���rW����f���%ޯ��1u$�&�����Q0�_H���X�C���S�&�7�Jpr�B O��1qVa�B$h�ʔo ���@0w�;~�{��>{����s\y�Ț�}��%�1�ж���Xb�t�pJ�]���X����4e�B; v���~���ؖ�+���A�ㅆ���\����uR�˻��Q��܁��2h�m�( (��[�8��ל`�}��C�5g|�4�UT��}�������_?�Up-ΛP;��r]u&^�_�I�D$<�g�b�.�OLZ�o8N$��~�P��f�?�S�=���Ģ�l�� ro�A)��ԟZU��I�9������+�����T59���F�`��^b��O�Ģ�=y\>棳Kn�҅���Al��zY*qÙ��q��~|s;��<�}k�|��l�'Z5�_P���"T��mʣ����&R�ʎu����)��w3�K~���X<9�^,pד�v3`����&ͽ^���ü䆬�� #���� X�ϊH@��L��r�9�i*O7My�B'y��lB:9���r%Wl̚��B� d?�9�+�Q�#�K����ױ.2!�Ԭ#H��-�3�F�٥�����Sk�!�/ge���G�'�}����*uݟvS~���J��s�n�d�}�Jt�=���R�e��l��DfY�����[W�0N@�fJ�ҔA(��_Huc�X5����[�?U�������c�$��-b��fKU�`T���m/)-��ND�J24�;�]Hh4m�\���}������9�\G�N���`��_-��Ə�dzR���7�k������
N�X�x6�����p�'F6�bG\��%����N�Q-�^H�2%:_%?	<��m�5�Љgq�Ý��!a�_t��m�h0�0�#���ۄMB9��tDp���ڠ���������K[ӥ@�{��D����W���2mǢiK�����v�L�RU������P�X�V�L�/}����Kp�*'�#���k3U�?!��q��!��x�S7�U�eǴ�B&�"��o���WWQ2���:U����{]	�F�<h%�u'�9ob�8��_�#sl`eP��#�w�K�t�Nl�h_�f�����qQQvc�;y��ݎ���n�y3e��ߤ}�:� ���W����[6�)K�)l���~V���o�;�Z\`�(Ԩ$�E���=��A<����m>�
|J�Ϫ�#��ɏ� z���C�jjf:k.`�U
��yKS{�n���c�|��%AƭEV�ۑe�~>L�De���&t�'���'�M�YCA֞Ϋ,¡�6atǶ�<G�	�IH�B}�_T�B�u�<4����1�������A�S�e�ofv���ba�e��Έ��x��0r
��+gf�8���{�|N���{݂31���)�`B��m4'3�dt\��O��`G�T����{m&��+�h)����;tK�q6dc(A-������5p���Mh�r/��$���+�rߪ�� ��N�������_1ZNZ���/Xā�n�����wg�����˲A����%�]X��\P��&�X�����l��F��6�ѣ�ϤtpTp��uτAt�.�+��8������ʾ��j���/�˕P��%oƭ��6Q[U��]}V��{κݨ&R�����4FS��=H�z�n���"6R'���U�E�*��J=*�����c�0�|�|Lߊ��}��v����0_�aX�V�L���.uK�$ǣ�o9xXlxVHYEB    a482     f40k篡���0���me��"��EY����x)�I"����.�����Q���E��#n}]zW�=�0jތ�ZX|�WMy��*G�<ϟ��%,�X�r�ɐt x���vX��;�1eOYP��;�#ZBz¡&�[�p���2p�Y�ԃ�:~ԴF���HKc�5U��`hy]So��9"�Ϛ���*�)~<�I�CXs�2̫��[k�Ƽ�LC��NN5��>_ɊD��M��N�*���[�V���A��R�:D��Z��սwhw�b!�ʝ:��j��Sݫ;��ƿ$��WO�\�� ���
��&%��f��Бe�-�h�n�� ���P��,���G|��f����z9@K�b4�[��$Ļ�:qQ�Hd$�)~0aJ��$N�]��o{�匃�Q�3����ڭ�e������(��2�5�SJ��.پ�d�ǪƎ���$�uG�3�:��8�R� j��B!۔�ּ���ԖC[rIo&ִuJ׭W�fD�V���:����N��+qĜ�9���C��b�M(F�2' {��~cL�
�ܗ�
ދR^. ү���)�ڰ�)��� n��O��l�)W^m �vyE ^=�gx��І����&����~�M�ݧe��2V9��rwC<�뮑\^�eJӡ�}[<��\�r׫E7AD�g�+qI�����Ɲ��/���
��P"+?RX�(��G�>�d���A	#�!�u�$���.���ю�݀�P�����X!��;Z�N���s���7�{���#���=9���*2$m0����[�ݬ��+y�P�0w��!K�]ޭ=�)`ǒ^�P2����>��Z���C�H�	�`����;�'��m�V��K����'���A��o<��~H�񯙐�w��
��&.�t��-�?��# Z��0�I�p����f����� ]>�i|g���[AT�ӣpދ2V�Ts�I!�ȅ������je`����O�	6��B.����4���ՠ����>p� G��1,/�{��iҘj��Î��^��X�u����zެu$�	k�FI�|&��B�� �����K���ŏ^z�^��\2���gA��+b�w�o���V�d؊<wm�ZP\|LF��"��ݧ�Yf|�k�����F��h���L�n���t�Vi�ծ�)Ԗ'���P�t}���1�E��?r7�� �Q�O�ZU���S)�qm�v�ů�9}�m��u(d6nu�����nkb8߳�CC�p����ë�Q����IQ!�(�m�:�Ǎ���)�K��N{27���� s,rb'g�y�I�f7�Ī*�U��$�Y� q�<�O�| � -�Is�73D�
*���X�B�}��Px������	�g��F荽��S�s����K�d5���}�<](��챹����1���(n��pHk*��-e���H�}���&)����Iu3GՓ�s�Ɵ"r���������ʩ=��$�R|+�)�s�����\3�mI���L��aٗ� #u��P��N��*�0y�b���`���k*�ok
7]��1s�.~����O*�*Y9�����0�ۄ�ˠ��i3��M�� �D{_ۂ��+l�Z�����B�m��s渔�$�T����hp�&���8�H=Ǖ&-�R��պ�z��������1�[��z9/c�M2eV��Xɖ��;0N�\�^�_E�A3ؘ	�Z$�?��4��߭M�jf�70N�o�!%�b�1��(����5��|�z��i�A�:�([)x�X����G��&D��	�m*@J�N�%m��_'�˦UM�y�k3B`����0��g�������s�NBv���*r���!�F��S���o�T&�L��%P݃�Oa������)!����P���OET��}L�{��ۦd� rؼ~R�W����NI�����ۈQ�򈊻�S"yL��������U�q�FU�}���F�|�lɘ�?��˰ڈF�S�u�k�{�A<A �À�J�A�����N�,y�)�|�ͮ�1�r}�oS��6ܨ�p'ߵ.�c_�:��\-Z8Ei^���ے־��u4&u�k����^�㲒�	��cB4����;<66��n��'7/�1�����5̍3
�\�ħ�fL������=�=�Jx�mZ��C��f�8����.7,L�������� %NZ�={����#
�g*�T�aFl�9C�m@�NJ絹LǮ�KeGA�Q8��0�F�Hc����.�uB����xkn��d������&����0�|m�L ��ls4f9e)4��f��?`��Є$�b��世b� �j9�3���ɖ�n�h�t��pŭ��eWo�� 㐱$���'��bM�6��1���,6�#5�f�lO�c/W+B�ťR�>�L��e��	�8��iz&�����H���3�/�`��ؽ�z�:���|��=�-2��|�>�~���4#�RSn��	�=L���5�#�r泣�МbH�����Xa�G��e��E!`s��K�猊�y�VZSA�E��}7�T�	v:B�o��?�d؞O��^ʙG%��'�x��TE:PF�g����Δ��p��%���c����7�`v<���-����Op{�|Q+ɫ��lou����(������Cw26c�=��Ӄ=9ޛQP)�o�� ����c�M�F�Ȣ?���J�U 9���r��$�'��V����(OFx��#��͉6���9&��+�o^���5��Zta� ƅ/��p3��_�X��'���S�5Z������+nYe��x>���?��ɚ�wol����)C	�1	���)R��U'
L9O���$ 3VJuwi�	P�E�<,� �&𵪻yMf�F>����c{ 5���{����~�ۄ�Ȕ���rK6���%�nBZT�O��)N�N�U.F�d �'���/�\�a��Y95lw��.Z�t!�q0�8��g-��N���E��ȣ�B(/�1\�[�I���˺K��d��^�/���?T �×��]F���S�<�!dFj�v�:_��`'�����Ik�*��ц���td�W��:/{6�#�E74 �R�
*{�֮Π��7vC�@FF!����w���`�ԋ�&�B�h�2Z=���S�Vn���,Z8�O�����| ���E�<b����0��;AJ*���?ؙ�c=8A���4�.D��2Mk���.f����Ͽ%maXȵ�tU,�������=���
�2��Ύً����n˧Q�b�>��fwHXhfդ���VO�E@֩w�w�FV¦�A��<y>��|N>��h��U�.m	�S��"آ���/D�a�ƭ$��H�mx?i����� ղ��M�'��W���֫{������+��Pd�o�{�)��IDI�'A��#/^-��/,h��Q�� �v�$�m�i{��}n]3B��Oya9��ӄ�Hu����'� �ܓ`:t�̫إt�W���	:_����Y�OT��4D����R�)�H-c�h��SYЕ)$�_�����E���������wb�q��bQѳY�)��>�n�0��)�qJխr,� Q�;�d�.z?\	�z�êG"�|#�|�1q�Q����@��BMd8Y1��g���JlA���wu7���9ڵ5m,E�8���*S|y=�sw6� ���~w��J�]ۿ\ۥ��e�,����΄�sJp3^RI��ަ|�� ?��4�!��~��d��<�IPgD�<_q�Z����� ��R׆K�Z�vv�?=)�> �e�a�p< 1Y�ba���Sܥ�t9�o���w��3SW̾3�C��x