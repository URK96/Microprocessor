XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����z���NS7�4�BGi�|<��u,�;KݓP�p�h}B�և"
��T��5������i�4���t�5�>�dx̩���:.�ے�q��;�ʹ��W�)<�m�w�M�~]��p�Z�"�P^���<~���c^�`��4iٺx{�Ⰵ����`��DBK��q�GM���KÝ_"�;�.�.2¦m��v��OS�9��y��n�f�� ���Q���z���_J}�Ho!�w�C<���K�r��-����l��3;�ֵ�z��t����(���Gk=��J��P�����d"J�/�(��YISZI���.�o��Q�n�@^�)lq�c��cY5r���<���Yeч�~�nJ�-j`�*ʢ:Uvs�Mq��*X
�*.k!�Fuv�5$�*C*�e�-7��~Q+��(����f����X6)#K{q��X7iik��H����{�3�s��n���f��fzD��;���5�� v̙pY��
�y��N��-�핡�S9�Q�9�N�>z�7oq��n�����~B�8ؗP������M�Z�`&7�� ��<\!b�a��Ko��1�}���"=���@fj�K2�L�u�[�8z�!���:�A���ǗZ��[��"�����V��3���ze����t�E�*(&��,K0��6�u��q��<���E�6�kv$�2(B�~��W�Ց4��ZDL
����eB��u�A�����c ��.�lzG�r!r:�=��M�����XlxVHYEB    166e     400�y��8��+���`�d���n	����^B.ŷ{�G�9�p;w
�8`{��D������j�)B�����#�jx%0˾D��1Z4�C@���:<��!��h�P6�.S�dL�$�	��}y̤͘"���3�']t+h�T��gE�H����ͨ/�Z��2��ܫ�4�ٚ�Н�j\�V���吮6����f�ȑq`�|-��zqݮ��T��w�}x��J��J1��kp��v+I̺*���5���{��E����:�%[�q���)C�U��"+��C]�2���{��ER�����mK�R�C�6s�����` ���*�OK� ��5g�Rwl��uŃ	�v�y?��)�����D���fߓ���g���w�9�r�`F�����ދ�|	��<�V�m��#5��p�^�A�1�`q|��>�H3�����8���R�����UB�4� 13H���^̙�P�`R����Ïsol"�U
�]��d����.��a`���b��RL��ci#s�k`ZB�� үJ4
O�t��fc^��2԰�w�_��HBx��K�R(��QZb�p�Ώ����p�,�}뇦QAA���>��a��R���E�$�n��>�xQrOD�	�ٷ�m3al�mfm�ſ��#���z[<`������  I�-�9�7lo�>	>��q�T�Ǚ���<2卄��*Yc��:�i?���f�O�p�ƊTE��	IQ�2Ӑ>�Wˮ^����}��!^T��tn��V,��9��\���]���i��� ��aU���R���w�|����1���&�=/�	�*X�0:����o����)��!,�X���U?J�Sh��f>,�0��t�o6��\�6`؃t
��i�Te�%Jҿ������^b9�KAvbQ��^!���% �w mX�8���^"��D��&	�و!�cM�q	��iP}~i�ǆ�I���O�҂��k�'1�0���=��F����N0����6;(