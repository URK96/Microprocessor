XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!�>؏ B�>?�~�m�~��Bb��������@��?E|�<mxc&�yz���U�y( �ӆ��+����Y)������ ��D��ۀ��(m8ڛI�r����Lﯔ,=M�4����ZR�%"z ����*I���G����0M8�T�lu�ql�qs{1�ּ�3{q�K Џq��
�2�l=�I,�/x�*�5(�$�z6+hsbY�{�z��*]��n?���'Z��ms��+�)�����U\������������}vh���Xʘ�~N����?�Ś;q�}P����j2��
���PeQ�~¹�����T��}�[�5 M��#��d>��Fi���I�Xy�A|�E�xZ_�6�4�Ú�o<(�ǩ��Cut�7�=��D�} �\�m�v�b1Ô�cC�PMI~�;�����b��� �Ql��8��%=�̙�7��K�V�������Z<B� ��R0>�pC�Ԝ?� L�2�Fr�!4�\�go
�^� �Ì�rs�U`�{��
����L���|0�������=Bp�ڡ�鋣9�$���po�9�S8��{Vl�េ	�!�i8���ً�NE9q��X�#����zN�5g<��R���@7ꈊT�i������qc�R?d%����=���2DOa!�Ԡ��1:�/R����;��my��]�Y��eK�ц��1[�~�w��N,b�?~�[^�%�������-H��uv3G=�I@󐎞��2�o�h�e�M��&1��^a�RXlxVHYEB    2d5f     800 � �!����Mu2�3<x�4c8$|�K���Co.�,Ȝ{���R&��,웯�cΨ�v=�/�p��3��BdW)���T��&>0�|�wM�ƿ�Yx ��6��3J�����^�5(T3]��|�,n�!<\f~���H���]M�ҙ�� �`N��oI.
9��������&_GkP�)�$�=�0.ʖJ:��5�%���i܋2~wRGg��P���%Y�Z��od)�~���R���`�p�s��M�iG� ��0 �p�h��^�\B7�8vr5yr1��8��:sC��
��{=VO�jr�'WĜn4�.�06�E��8y���_�P'�+I�ĺ�1�b���%wd,}Ϩ_�މ�dB��`�~�>;tL�Y(���1�!�#��Ƀ���CR)5��'�o�?�\�X�t'�.�U�������;TG~5톖�C��V���{Y�w��.oy`���A��*���T��{s���ƾ��`U�k��0�;�  v?N�Q����H	�z���g�zT�'�t�=���|�/+��Ɋ��{2Q�P�ӋZ�H�GCw[��XH�4q�/MG;ǿ*N��ߵO�O8�� ����f��>J0p�*�bR�+\:��F��;`�����C�)�4��[���Js�-
t��Xս�xt�G
M�Zj�ҡෝ>�4���R7���KV�0����P�͠!��>��T�.�~!=
Z�x�'�v"��֤�%F<��J�B3���=���U�V�oUD=���,b�1��Ĳ�<�ƙ�5���e>�QVK]`ᴡ8��V�>ZL��N���ŢΩgy��]�����㠕O{S斓��u�H��E1�_�_��+xi�^�C�>���8+A���i�3�ʎk��vC�ڼ�v�'�!��Mu^O��g"	������b#Nʧ�S2'J�V�C�h$&�3tMF����α=���.N E;.�q���4�"G�j�����:� L>���Zh�#��Eѓ�=��5���I1#�(	K�������a4��&��'�浗��&�0���,�gb�W"�ˎ�&�Y�{|�KvRXs��}�x�=��q�w��wT�g$�Ӣ�� �F�z����f۲V��P|�I�P[8��Gn�-̴����h�Ym�^���Љ���}~�<���;��.kz����?=��$�C�."�V�<�\"��N�qc�R�V�����^k���-��a(�5�C�-a�<\F�ѫ�^���� ���Vo�`�"��̡K�C� ��4���D�ҵ_&4c41]�8��঎ϡim5f2��7����K�N�hJ�\Fc:�cCj7��;����������E��uk�O5��@G���h� {ͣ��F��R��!C�xU�����f�;����L�hܠ�3���(H�rz�8i��2�9T��(��"�*+�qSa��D�W��u3�0,	�����t���#��Z}�,�X@�{��p�{CW\��7�E'��Ў��o�F�-�5�g��WYҢ��V���]}o#��
����Q�G���$�O^�Ʀ��]3T�Q��2埔�wA�/Ƽ�%�p�^B��jR�ǸEL�~g�10�3+Nɣر6�CX)�,E{kP��v�v=��-M�K}ױ��x
p��g�q�fۢY�/�cL��7:�|�
B��1o?8T�1k���e�b�������YmgH�S#�j��}�T�6��
y|�=�7����e�t��͍W���R_@%i>p�����j��Eal��I���R�gͣm�׎�Ǯyx�޿+��rAK�7�ʆ7�ף7�i��lx�j3��?���h��*P�!5V�����`퉤�Q~&r��"��2w�n ��?�*\��|��� ˝��z7Cb<D}to3�·Ur���Li�o���q*\����|�?m��{�Cd�ݲ�2�D5聛
6Qc})�i�r��<"�c���q7&�	��`Y��{f�v)5fI��v��[�o��#UV"�X9��u�� Ӄh4�