XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���7��nu�����v�#�We�^�ۢl��Ե�v�:S��t���.7["��ҕ[�@>|	w�PhSߡ|E����c�N�ԻН����>��',�c��O��	'������+�Ǫ��`	�{5Q� �����v���ؙ%�MK�g��&h��VU�-�j>�4[��>��J�D����LΑ};��\�Ci�C~�ݼ�P}�=]D���9�h� m��i����{wTSyZZ0D&�DI��]N�=~�X�-6��
R4;f��ɘ��w��.�6v�:���
&����5�a��?9>n�$��!�`[K��Xu��Wв=�i���:ĖP�f�
t�ؔ#�ZE���	���g��#!%*g&_�Ó��$7$��\eW|6p���≀L��
g��ƪ3"D$@�:�V���j�tt��v뱱�x�u��È/>�F���Ug��>YxzwE]�y	�/!(3�.;|�e����$�C;RTXZ񢃜$���9�I��g�����MY(��(��#(`K����{��Q#��$���ՈO&[�o��.Q9lQ���S*�S�*
N���L�;QQ���?�̓���4�[�޹+UO욗�� �U���;ϹJ1��1��%?aw�K�]�Ԗ$����k5�j�aU$3A��F�l$�Z�̌��}�Ӓ	���J_��u@��Y9��}ſ�DgJ½�a�Gm-(�j ����ºOK+-�=:�+�R�XąË����_^,d��Ƒ�"��Hbd��XlxVHYEB     705     250�L������y� .�z�釩$G@��V�>À�q&�,�l(9-C�eh1��ex��@p�����f�n�ĭ�,²�n���{֭cP�L���c�=�@3�p@��\H/�\n�}t�̫`Jl���]ֹd�k"S39��r�Ů\Y�*D�+- �f�9.���Qh�c6L�{�IG��|:a.�Y-65j�Z��b�gH��IDr�X��������?k_�e]�����|�m��כ���*����C�&�.���Aed��ɯhz�c|�?7�1"�fh恜�������$�G����z��$��X�;���y�,&h�0����?���#��q�M����p�K�����x�� ���Z*��-Y]����J���(����c�5~߀��0�N�b&����v��"�;��*x4���;Dtڂ��|@����*��B���	��2���O��Jm��^�?^�h~y^�Bj\�0	0����H�n���\\C��v��-۬EH�����fe��N"�Fr-j-�o8��,WB�P�[+�#��J�3�\P�d���ͧ0��'NX�;=����ܲaQ.��t��WA