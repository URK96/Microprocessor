XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T[.c���?l��h9w�a����4�'<�=����Hbu�h�S��bDS_��C��3�H�
(����N�&����@��?zhV��.�Q���}�L�]-���=�XpE��0�Q�l�ܸ}W=�j-�X��W�k�rG�l���w��~��T2lv��IsYJ�E���L66�J_ݷ��4��-b����)���J�P�lg���M\�.�9��XQD�e˱ab1&(����-�w4ȝ*�:����)sɱ�kũ���+8��>�'����	;dW�ޙ���0�O.�:��pU�|�� �o_�nvx�	n�1����œ�՗s�*܎�%�樦tkhνT�&���nv����Q�k!�Ơv��i}���_
���ɦlҀ��2�ƃ��}��P��(��
;�~��oOhf�L�j-p
x�qD
�02�X�"c1xd��Ǥ*�I#��
H��z3g�سÓ�&�K�~�7Z1���>�k��c�bkR��lϥ\Z��� U@�-��$v-wi�<�}��񋀃@Y�}\)"n��q�Sj���QVl�r�8R���`�.X�<��]�מM\�\0"6�S��N*�iGD���V� G���ƞ����ޝ�c�0wiĻ�e8���ߑ�tP��Ltq@u��-Be�4��0�]���ȬĒЬqK#�b���1��kr��>��� �O�Q1�)~�y�p����8��Y�a�۹�n�R �Fސ�N�}D���n����ޒ���/ܴ��$\�~O�O�'`�UXlxVHYEB    225f     610�]��%.[I�Zu���S_��	lI�j��>�-��t� ,�{�pQC�w/�:�a��>e��]IuT�/D��eAUn=�M�uT�_Q����O��= ��d�!oSo+ו��7�t��C+(#o�a��5_� �s�T�����,��xQ@8�p�iG���6b�q]7}�B��/5�'���淣qd�A���cm�����s�:"��V�B^�ڐ�w���������?cM�=��f�� � ���Z�:[ƽ2����[NS�2Ө�N�U߭J�U��Ȅ�n�����`��`Tz�ƾt�D�+���J짃� ��dp~�`�3�:t�M�Ds��sK�q�~ ��B��=Tw�#�I�*���ʽԆQ-�(����v��;)���q�i���h'q>Z��eH�������?b.iz0�w�v"�5�\Ci�D�}���K��L�~@V���\@�I��rRTkC���߯�(A�"��b�j���4���̐�6t�فƍ&���Y����<�N�b���{dE�n�Q1�Ю�*"B0���70Z��Z|nw�=4�۾�낔�l�^>��G��+^IFc�n`��F��#±�V�[�d������V��S6�u(@K8��7j���1S�Kh�I�[�(�Y����`]I��`�hIG���1e
nC�J�GYww��PJ����uGW�F�ǈ��D�����C�ф|?dMIs��3?�R
eQ��ܲ��8��t��2��XX����ԇ��EZ;!Y��B�5�S0*���2�U�D�7]���#\���Ο�?O�;������O�������z��rO�w�s|�hS��f��6�Ժ~�W��7�:]B�u�90�AG����mJ'���;�l4S�U5lI]�-a/����ZT�"���G��lV��=cZmMD�BiB�P]�u#��(5$j3�V��U����V�q�D{��$)x�WX ��X����������=���q�y��)'C� �_V~�bcд�j!C�$����ml@ߪ�;�I�#1���N�1�wB\+T���_�>��6���0��:�c�8�7N���b��2�y�3��?d�;T��bϭ�����1{�s�'�ѾL+ � $�2��ŨX
�7��J6?>��lĄ��Zo�M^+'��R��dW��|pZ���{�8�ԔK���!�7�" �(�{0����s\xً�!/�K���n3d���-*�<�%�n��u!'? ��O��Ӽ���5����Y��o���vk�r-�ah�Fʺ+kYĊU���~���GrzU�w��[������� ��,�A}(N9\����Պ3�w?iʏU%	�����ogqVGS.tM��L� �T�j��R�b��E�x`=nS�
�5GW�ݩ*����(v=��xgu�71��54۠*��r�uR��1�;��Ш6��O�2��CG����'T�f�����?������[���+0ovmLb��j;�����s���5��9�Qt��mpk�>Xj�@�V��$���