XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����&���NJw $#$��hL�Rh- ��s������{GD�m�T���Wk�m٥�d����m�ۗT��9�콝!Jյ[!%�x�N�IN��� -�:�uH"�EV��F�~����G��Z����t$��`�i�~Ť������3U�(��'p�nm�r�S�A��?���C�P��8�lD�D��t��?:���GQ᧝�l�o�oLU��<��F��%(�Q��nV���m&���e�32rAcP�07��1I��5���j�WX��ؾ�ɐ�{�a���x·�)��X����镓��xp9����G� �W!�v�'�e_��J��b��T� �ҿߣ.��w@�f� bpm���L���2�r׍�~��4"��OQ���[��aq���X+��C?Q#���z��������oě��֧�y�������&�w<�:�Iȱ�e�8BBNJeb���Cz����5u�v5�v󍺕2���v\f7�IJ�f�c�����`[q��,f�HO@
ϑ��4�	w���LJ+U�v��w{�7�NP�Y�=�<cP�P]앏�K��>˭=J��Y�����՞�k�K�-����#!d*(}�o�T���Bڅ%t��&�����k�w_֕��M�۶bH����cy��$k.�Q�;��ƽY ֒ml������U���4i�*���+_IRKlG���t��)L��i��,�o�z�H@P�x���#�I�+�����^�D�ps�Ƈ�DЎA%	 c�]�ڪB�#XlxVHYEB    38f0     d30U�ϤA��Mv:������Ua=����WE!ӟ�����n?�8��R?�ڀ�����y`a����¸�o�������,�ҰgQ�*����'ѩ�"\t�N��w%9+u�g' W��[kZ��C)d�C<H����C�iZB2��J,�&�m����1D�k{9�U/m啺��0���P�>����'?3����,���g�T3�+��j��d�n�]��at��s����g.��.����	��ɠf��ͥ����0X��t��[�q`��Ϻ߰��"�)�q{g@c�*�f�J�p8��Z��S�H���&���8�qVQ���c� �S�� �d��kE����	�ը+��~�16�z����q�[�iv.��%I�T2�Ť�!�^tA����e�>��G�'8�s���g�q�8��(ŋc���3�Nh�y�q^Qjq�z���N Ƣ0P�/`����^LP�8���A$ͼ붅X�oA#�5� �0O��b�I+oT5��Ò���417�w��>)�7�IΧ��)Eb�V
˪��o�:E�������?x��1S_p���DŻ��u�P��sێ�6����	���0�3;7�19C��a��.B���|M���vN��N*ȟ��@ȇ��$:/Q���\96���í�"#jr�҅�|rS�o��"�r��y�p�1E�>ʽɏp�{�/�X�W~��XMֈ��yE�nA��x��}����\�jW�)B���ao�:a4b旭�����%��0�	i9G��;!B*7)E7�q�5��6'�['�1�:��B���F$� ��9��2
�G3��%X�'�1�d�*F��Y�v�bk���o��Jq�
���ڐ��/b�i��v�v�*������}�]ڶ����䇲s
m�
��SZZ�H<�k�C�T5���M
�o+ ��'{���;�|'��t�{�U�c�wr�/l��d��^Sh!G��X��/0�����	܌>_���D�%���Hz��{�6��p�PZ���%E�2{��U*h��ҕ+x�hP��XQ
�Ѓ��!
X�>�@2 �Iv��x�>[��֌�?�C�L��:�t<rH?�H8M}���^�u<�����.��,җ�3�* ��U�"#T��-{��U|���;M�b�����]�+Y��(X���*�R�sQ�����Z���	�G�r&��S�e�!/�-N�Ι��'�u���}����p:L���#������m��ٗ��Mr��5*�) �D�ؒHS�ǛW�:�%~eB��$���0��Vf��Bd�j���l�a%/�G?�|2Yع����I�G�7�v�{�)�a{T��#�UIb��/���"᪜<L0��t��!/�9��g�4���eM��xE�.ڵ��l�_Hk̒G���t�O��Ư�ը6d�|�N�Ȱ|Ѽr'�xu�����Y���ﴣDBn�����m3�N<,(��F�ɰ%-ݟ��� Lԑx!.���P4�$��~Z���"_W�}caF����͸~�+(w�-	N7Z�D;@Y4�����1���	c������GN���.,%8_U p-~�7ڦ�ҸV��o=Ԗ�ב�ǿ���Ձ��ʑ,f�� ��C�������Z%��Z��r���\��J��Rn�>v��FIIG��5�Z��>�w�ꅻYgDqo���$��l���{0����7�u30��V3�������g:R�K�T��ۜ/ت�o����[I����L.<-�*M��-����$�i�+@B�7���N��uT����Y$���n@����#��=֗�;���h��%L�Ht*[&�:\h���9#�@��!�����੶cϝ6a�7?s��@"3w�@�O�	��V��R||��Ţ�c���Y�/��҈��_�=S���a_$I�d��Y�I��R$���D�v⃓|�Xh��x�L�H�u�eb�5�� sns{	�-�S�g�y�EIY�G6d�iB����!�,OQ�����k��={�P	^�3W	��%d����w#���?6����V^qs94쓙G����^m1�[+�<��(�7��U�_��«�A�U��=$��f^@}e��]���,����K.��.����;��/�0Y����1�ۺui���n{E	+xUG�3�N<+��@hY���j�d����ӖbjF�-�.���-�n\�Lja)���R���(��-e�+_��L�7#ֲ���w\p	���"Ei�a�ǩ��O�+�o4AkW	����k�[�j��nAV��[��+�Tkɕn�$v#~GmH����f�vhI/uQ~W�����S6�Ēٿ�	-<8��7o���d��%�]P�p��7���bx�xb�ƹe^}�F����l��IW�0��bRγ(�@S*B;�m�-�l�b����7ϴ�u���e4]�T7Y/�W��# ̤j��&Ѫh=����`�1&M��<�Oe�<�[{<L@Sp��9��� ���Y-h�*�P
o��Z;��AMt*�S?�h�`\`�4h4�#+����$�(�)RT�n�?D}x�-Ye�����Eʅwr�oCZ���%�ê+T��gŚ�d�pl�<�b$��0�N	����gT,�4.�$o6��9���*}>i,���G�L`��>$<��*2���U�5�=؜9�:�@���{��e����7�D���X�
���}h�-�!_(��d-��@�OI�"��h����nt����u^jJ����%63��}�q� \�y��C3����,*,;R�a!��	�d5==H�Eh2t֔/:���E��$)�*�Ų*P))g�C�8������㓫�����,��{m��~�b��ԍ�Tc����3� u�[8�W��S�}آ���M���G'����Y)ME�	���>�R�b�Ԕ���<hB�Oe��,��ȃ���QF��n~Ѕ�#��KV�0�DF�qiZ>@E�����զk�����ĩ(�
%E�����W6;^��"%5�f~Υ�2w��"(�ٻ@�^���T)��K������� 4��oE��� �����"˂��r��٫`�x�QrH�b���"0�>��b1lb�L��MAj���~A \Ju�[ܥ�,H��)�-b��)|�u�x ��2�N�,���0����d�?�$!YRB�����T��e�g�n�L�ͺl�}fXĎ_��6'/Aq!��Kn`�q�O8���?bkk2���#����޼�%����& t��Q�C��c�g�JB,��֘x������
{�g��ڱ�����R?�_9���+�zo(��Y��K�e�M�ô���e�OM���]G��m=.�#��