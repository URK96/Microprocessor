XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E����SQ���i�=g����x�0������ ��S��y�A�f�1���ѥ���5�Н:�@B�n���X��"��1��/��02C��~����.���!���)��9?sW��5������*�L���l3`��mk:��>��ӜT��J�;K..�.��Pj>ד�Y�Oߒ�ZU��^4[��~'^�p��ЃL���bQ�d�Y�������{E���d�bv%v2���fz��@���!wyA'����������O�����Ry6��>�[�i�Tfs��~p������$�O��'�2�ty����{��kC.�3�����+��x�7�6�YD�X�KG]� �J�#�s�0��`�lG�ħ��3W�wcH�|9��Ԛs~��C~@fM�X{�� ���|}�u���?�'7�����K������S=_{Ѯ�IZWv(�$E�D�$�k�fm��?�Sb�xaM�������b��z	k���Ҡ��ځ$c��rRd��:6�<��!!��(�d��1O� �G]mT�ԓ{���v>�*��p	
��|����mV"jau(_����B�V�=���S�s����2�{��(���r�>r����*�V�̗�{;�� &f��-�p��O-
0����X��fR?]�1=9�~�oeG(�)(M,��&�Kqu�qM���gN�k�&�M�Ѥb������2�7��yc�ᢙ����K�{U}B��j��]Q[QXlxVHYEB    6fc6     c30�l���2��s_'�V�:����l�H����޲�`j00��m�+���f8�ӿ[6�d��P�mc
�V4��zYq7S�Ig�ynX���()<���8��ËSۙ�ơ�@Ġ��O�u���P�I%����Tګ���N0�D�.�p	�3(��1ۏ:���Z�W�Y�$x�ͮI"R�+����ĞV�����o����m�m�B����"���+�SR\�� ��q��8@
���!�o��K(��;rLq~�NZ�x��r$,BgyvD�ۮ I��9o}��˥��"�±fd%��l~�S[���?�O����� �Э�Z����d�top�mC����;�2�=�
��Tp5�}�dT_)� J�5#��� Rޤ,g�Պ�omr	(*R�ʯ�s�;�ܲn��T�p���#^�d@�-��8?տ�`4s$�3o��|� `�ԅ�E��def)6�8_o[���l��!H�����2_��@e�Nj+�l���oU�QsdҜ�z�8�X�� ڤ��ӔM
X�,��5�E�l�+]��M8e�y�����F*z*0�}8�f��z�ޠa�<���xL��5k`%�or���nMq�$Qx�6�rP>���ײ�wsS�jC�AY����h��f�!�\���$��G뿅�Ţ�


yu���U����G����Wo�/�YĜK ���B{��z�rL��՝o@�->H�����*@��O��u�Ky�h�N3柉R���iT���"M�]S�	�~��C[b3�\ǣVӱ��maX�j�������Q
��&l����8P�ަf�]ۿ����H��-�����c��[���P��V,�:��ץ���h��<��K~؁Sr���k�r	�`�k>G�r܋ma���q�煘�$��ޮ*��[���O�}-!���ThQ�e��rԒ���|i�>h���v����Y#��!BeS�\-ө���!��7�����u�E�|up- �$aF�!��
~e��/獂�H��ȋ���a��A}(����u����d��!�ng}lȜ˜>3��a��9u���1jO��gܮ
>o%���;J��9ME}#h�A8��=�0�S����St�IPj=b���I�=L�+��xӞ�.*��#��Qv��P@�q&n���Sr��G��N䛅E7t��K���� j0-\{m�����%������Lk�.KD�|�)��&�Q���f��u"2�K��ڄ��c/��|�S�#d��β���
�dj��D���:�W�������֝�A	/�i��t�Y�R"�"}$R�Ӆ��-9b[h?o�H%�Mp̞`TND��~��)|�7- �.8˱�$�԰A6L�N�H���<������-%��1�qwT����/��=%�/�	����j�D���������\�E?�An�6�ݔ?x�����L�R��3�z��o؟��gW_32j�^��'��I@�k����T�e��5�Ls���4��w��<>"r��K�8�B�ˌ��h㇝�;�G��
�X*��	R���#���ת`'x{���t�O���H����4���,[�g(�Pc���4�]>�ƪ�B�%W2�%x�D�a]HH��j��D�)%�������	K�S͹��D�Ĵ���L��㼩�N��/�VS�;@pj�78KU{���C��S��ɐj��ρ(������F�3�sd����}�˝��k�	�J�ϭ�w~���V�(�y^�m+%P~I�qM��)��)9�0v	�%.w���c�Ff�*tRԒEUWb��_�]��˷d@���ʮMu�էh�i�u�WA�I�Ս�݇����HTjo���Qn��r�o���2	ڭ����(�h��р8@��p�a�E������Z�8�sa�$�n䙗��+�3���i�3��eHN~��7�BؽA��8�()y�0i2<Γ]x��׃��p�o�zɬ�ZV>�DY�u����B��S�B�c�����A9��6�<����:[�,��[2��مk�.-\��U����z�R������r|pb,=�op���Hz�E�W�OB�p�)�SVpT�R���)7w_ K��9��ukrJ���)��L�1�|�,���I-݌���t���fB�
eR�[hƆ���Se�;�\GEvk�j� ���ɢ�U_bo���!	C�����7/:%x���\�=����^�_�go�Wd8������E��g�6K���fq4,�t���.<Zx�R͞.�Uk�a��"g���maz]��D M��S5�xUM��Z�#_7�!��	�o$a�����3r��K�DKV������7$���It���M�	h���,m,��:��L^_���v9�b}��<�*�}�'NF�d�jq49���z�ٞ��.����*�[���#X�`���x��\4�I~��ܴ��v��y��yIꌷ��$�K��6�3����Zϊ/���Mt>/�F�i��늴�F\>u���A��V0�;5Ϗ�)}|P-N]������<�cQ�$�]��ى�	l�Ő��^l�S���F[Ѓ|���f5�H&leN�����ܔZ̈́$��s��+E1�Y���$��u�{^_fc�r8�HT��~�������M�7�qX���GM�W�g)��Q��t<���W_�"�9�vr��	�;��#�?=,h/�bM{τ(�����94�x
ӑs�_�rcrB�]� "t��b�+ϥ�:�v�T�+TJR��$��Yk�v�δ��H�hTF��iS��/���5��FW(���\�"}��^;ѩ+�{��eC�߸(j�W�ݭJ&��Ph��8	p�2���qì�1�L'��C���7,���R����X0��q��"B�Y�nK�E ;�Ň�ե �.�D�f��(n]���A�֍0 I��D8B�ނ-�����k�/�e��雒ԴiNߣo?��^QT'b�i��Y2�ʇ�uZT����o�|?9�]%�q����ȹ���A�%T��lF,���~ꆎhd�K�r�W�rQ���H5.ș�j�Q��z =�� R�>�8���2{�J�ߜv�qE	�3�d���1�6A�oMb�