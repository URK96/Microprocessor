XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X��]KK��������%%���eH2�љ�b�NY�P��UG�R�"���BE� в��s��|�î���(O�~�7�r�����\ܨ�<W�I�r�Q�
��W=	�\�܀��g�����#����w��N`p�Z�	&LeOj�c��3�UZ� ���bY��rF8YN���)a�=� e''+}E#L�Z�L����[��TF�����M�M.�ʄv<�t��o�6�fj;�_�?�n�m�VA@[�&#4z����й81R��!����Ӿǰ`v/p�E�@�Y�;����`���. G�������8����Ea��Ł��
"�U�>e�4����0rĨ�;g��l�M���.����N�:���܉��,~΀
ng/�E#gd�baJ1�Me5���^3M?#��w�Ϧ#`|�z�a���WU��o�L z��h�r$h�X�g����q���ޓKD�-`
Â�6� �b"q�!i�/Л�K���P����e�H�h`f�@�*8���Y�X�"��ٽ�i�����R���tG�T6))C3`a�L3��ɜu߬���]����n�%�k�T^r�f^J�_I
����t#���#Rν��.�Gʶp@�o!V��ڪ�}���d�\#��W��ydnF@� A���k��u#�J��$kȏ��Z�?�_�=���ql�ȣ
���ǟ�z�&!XV��xT�x��V�`2t�Z����=��TTc����!4���o�#�.^��(T�6T]l�^�f%<D,XlxVHYEB    41c2     c40��r[{�tu|�f-�蒪���	*.��D���Npv1�_x2YK��ߚ�S5�8ۀr>���R��Zr�?a(����~�/ܸr1gDe��P����G3����B̭X�/�l��t_�vωSh{����=�H��Պ�҈�-rJUa��
Y�(�x��p&�@��y��+aX��
�a��x+R���]���UTt%L��ݬ�~�1���`vU��$kĜA���5-���O�bi��px�+�?`_a)�_  �2�x�{��
���#G�"�����жp=d!�r���L��,E���O�m���C*�ߔpfy�d�=�ߗ��QI
`F��R.zQ�c^2H{[h��Y����.�*`M�\A�7{��n͋�;���JM�kǺv��T�	`�B\�W�M�k�vB*cLb%��~$Y�Vc���do
����A:~T�(���x�����C�X��_����ӟ�D�_w?��$<jy�n ����U�f]��H�AⒻk��:V��]r���C]�N���N�u�Nk�gJ��bІ�������㆔��4 ���J�Z|�A��yy�(��3�{�V�z_���-�t��BW��ȿ����<���J�f4�
v?{uU��"�v���:�����{��Ԥ�z��(����S�<	��˷{�)Q��J�'Յ&��5��a�#��^:��Z(�#vz�km
��s��`"ۺ{r�eh�[�'�?�D^���I�����Y`g�{�r)V��~?��)��?��D�����g��!p���o:��x�g�ؾ�I���%]��x̹E�ｯQu�����x��.�U~�6�_�a���!��U��	��B1!����$+�CR��(��k�I����Mbw�����[���\^�����ǆ�v�H�i�r�u����t�F]v0���X��=��Q�����
>���㼿a��)�*��<S���+u�?�&�z�pz�jtH����TS��{)T�摄9�((Q����5h%7Xj�n��	��P+�ܡ���Ӱ?��6�f�E�&�<"��8��@Ǝ����cJ��y�p�������	�� �ȰQ#� �X������e��0rR8Yd�`[��Zgھ[�MXF[�O�-H�XSWN	R��?"�'���wHۼ�WBI�ER�E~nȬy#,�mIQ�J�I��A�y�CG�c~�(�g�v�����[�R�yZ�Fk4�9ɛ�N���F��ʬf<�!�]�O�HmR�k9��a8�=.����P��W�G.^��l֟���u`�mC�q�PuX�V�������Xa~����W��i�&-��t���x�¯�pzx_��2��5�1}��ly�Z�?P�cmN�Cq>`�e?�.hٹ�6�!¹U+x]�Uk2��dE�A��:�b*��������6	�h�Ƶ��+9@c�H��)�������Dk�"�=���%���g�ΛHe�IJ��.a����4�����L{�k��w/�8���>Wz�J2�i�RT�\������ 5�,pY{(1K�]t�d�����=T�)Y�h�*���B|�ԉ�Y�# 4|>9����bYP�s��=c,�u���|���7q�1�����\~�H����(�V2����^�WR�Y�����(`��jC����elR�%C8��qlu���K�VW}�0�-Go8'^�'��d~�R�Ώ-��~gwe�b��?u�3hʎ��m\vFm�п9&H,�1/��FFw�wP~/�A�^y ���3C0@��bEv�$�'����e�3B)V[��V���{�Њ	yw��A��$���i���� l�$�� �Į����P�O[h��sK���puV~ �Gwǎ
�_k$tB)�;u&��-{M�ՠ=��&���:i�K�=,���C=����q�I29r���$PQ�x\Xմ�熱����k<�L�;f�~
�ˎ`�-��I�y�+@H��q?� �~ξ�T 0�'df�y��k���~#�ڐs.�q/�<��;�r)2��B�[�9��@o�~�'�����g��j@���� ���"�NgeF���K�(f+v����:L�HUfL���Q?��*��9z�s��:Lfo�Yd��1��9�܊��۹L�X߬��P%��z��
�_�}�c��$�%�x)�̠_�%�&-�8	:P�fQ���R*
5�Y�
���4�e��~��}�,��>�h�����\Ӿ]8�T�	��A�;�sk�V8���TѤ���ڰQ�B}��&x�۞D@R8ķ��d��B�#�).ꔾ���+%�NA���^O��ls.�~b0U?�o#�'��)���j;}�iÅl<��0
�y�S�� �\�@|��i��T@������]������Ec�r��hM�bp�BL�����
�^�5�Ul�d�er��X���i�.3k�=���6V�0��'I�1��pY�@� ��鍗�V����>�a4m�5� ��¬�pu��p��p��F�Kv!�	>�}�.����B���;h�@W1����@+�By� k�r�_�2�֪���R�̪m��=��e�����m&D��0﷈��-r˷�	�<I�����T�.Ѝ�2���S���u��֐��u1���#{�i�,Fk�>��@�	βl#�j�sٲ����_�<����m a�F*A�9�iLF��=N�3^H
���#���Ɯ�=�9�i�a��p�-�p�I�65�8	��d� 6[E�x0>^)�y
�F�h	$տ�-�X�� r��˧�bq|nJ�F0�DER���$Ҳ,��ˉ=��P0�(��.�þ��콏�yn}˨���{��s#�t��9<�|t�B��V_��V1��p��$�yƗ�C�9>7�?�H�r��i<�����W�H�\H<���s3m�2�'3!��a��{E�q$�z��|_W�//ɣ���@.��Y�	��*��pUE��e�w�����U��5CXݐ/���>��tӨ�TT{BF�Z��|����^��j���ݬ.�'��y�/�8��F>�7����fT�i�����$3�3�c���g�T��f�`��K鳟�-.f��v���}9�