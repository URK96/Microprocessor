XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��? j7z`L�DGZ���09��.�JeP��ɥU����-��8�1��8A.V�����x��{�k��k�EO��#��w�	�&��.ͪ�j_j��g�}��~	�3�������A�>��o�<嶴���[��SDA�S{ǵ��i�*�z�:J�\�{�j�)�W'���<�V���0���Qj-T݇%�q��X[ #L�\=&��'�1\�)M�H�5d��a�f���pu�
�]aK�[�k��N��V#T8�j��H��!<����DԨ]�٦w��p�-,���߸FJ��H!���Lc{��ݻ~9?S���s���^�D}���ߒV�QX�T��/8��گ`n�''k�T�]��mԬB�iT/��1����a҃�b
����'�\�c���.O�i{.%p��R�)@2�%p�"1k�e���P��N���mä���	p����Q�Lg#J��~*�v�(��[�*�:����ZD#�*|�=��FL����kp]mB��KI0ہ=�ۣ���0z�5�eP�i���ut�~;�-}O���h	�u%S�#h�x^�'y^��W�zP��sM��vlp�x*��'�+X%]��}�a�ݸ�#��Q��p�z��4�l����>�~:n��T�S}�7�j���Y\��c�sF��Sݑ��ӣ�������c Q��e���.$z���F��W�B~���+�.Xʿ�{�m�T(�}`"%��Ș=7g����V��	C����D���*黹��C�XlxVHYEB    41c2     c40*vQ��e"7�%�wj(Nk#E�Wͭ���!@L��p\aA�xyg0�u���ܕ������L[���A?L�T]���du����2�⧃�]"��k�m�����J���B}�wq�Q��*�S��h�a�{���`0Z9�5h�i��_�� ���Y�@�rͲ�^u�@H^��^���c���74����ӂ����1�5f����_��%$ʅ��^�����W7�j^v�J��{F@c:���H
P*�m��إ`Y�B}J�3".��(�56RF~U���og�Ώ�{�elw��2l�k/�ɉ;m� �w�`���8��G��k}o;�R.�/+^Nt�2��Q�9QO-����� G�oCR�/rmoU(1=������~���@	��'Pݵ%�8��j�R�KKi*�m&�Geey��B~�ٌ�|�W~�%�<7��4
J÷�V�J�a��׽c�oiFp���r����s��-n��J�L	��� !O4R�y6�C��`����k�b4b�����$�%��@�X�_��]��?�Q�&��7�.mȝ_[^V1���II<rf|{U��Řg��Jl	���;����H,� �EF�n&f�sj�+���w�-x:�U���)����`��k��Q�(�0}�I�,r {�bjX�1%�(�(��Z?����J����e�NPy�a�}`��Q �b`c�I&��/ʃ� R����7W�'�������!!b�R)YNm����ɕ|�*i��!F�
��'��ʅ%�楝�@�7�K�O�m ��SD&���ŲVu���ExΎY�c��h耬p����@�[M���;iq�>�x�?���^M @��ހj�;y��jy�M�xv���<����_kL���8�F"��c�c8�i�p��*��N��˫f�_��ܨx�ǲ90���V^��Wu���V!*FYIi�&߰�h��i��'e:����
��,��%����� �2��{j�e��+��%�ťg�XR��+2���p�9F�@�ۊIm~C����%�
��.�%�{�K�&�24�vvx�-c�kN	E�/7�_#��:SW[�u)J��IA�٬�E(��ho	���MLR猹Y�>o�űS�sJ��L����!�O}��<��JD����jb`���z(�G�B�q:{)q�g G�kɐ��L��t%I�֌W/ns}��3��R��u��8ę˱&�s��
�F���>�w�}�+^x�z-�)�'��w
�������9kx� �ZQq��b �֡O1<����P�EpT��wq�mFk�<��گ��_XE������y��7�(�5\70��:~J��31R�\vM�$�dwM�o=�S�Y�{�.�@�#�T�L�l���Xoֻ�v��e�EMiZ�0q ��m��7e���OK�ڦ������ឱ��EP�L<c(��#��Nh�)�>Y�3���0P��L/y�,���Or��;��~���"D��Xn0�� ;&?�	�����O*������0��5�Շ�Y����)K�������w�Q�{Z��N���@3 ^������/v��~�'Pӻ��n��Eԯ����,$Y1`��8%i��|�sб�Zc��2��*p����H�#Vc��.^'$HJ+�A˿�u�:���R��^	AW*n<��U��iC��
�W�3
�����R���T̊(�� ���9Ac�H�<���>�-]�n�h��m�g�e08Fx=�L��Sq�\@z��І�2��� /��.7�(UB��/��o+Ǆ�NV�т3sH3ZF)���ֽ�j#�������֨%��x�~S\������I�jZ������]H���r� ]�(��ʗO�+�Ir}�u�{Di sJ�^�KHi���9a����Ak��H��� TWCo��̒�3|h�H�HJ��_���ŀ$�8l��%~���Yq5&�>e�BE�Z���-Ȣ6��L�'�o���8��bY�&��DAo����s�-���Y����b}�q��j�M�e�,�"�([M.��M�Ϣ����Q��L�`��*z+L�����#��*���|5ҏo��ف.�`7M���B8�6xsZ�g��S���ׯ{>�A�86�<���^33�k�����YC�'��r�� ($q�:���KG��3�f�;?b�V��,DZ�������Za�m������Y{c��_5��.v}�a.$=D��e��C�i�>k���0Oy^x�$������Z<�{��\ʸ�{�,����V�M�T��3��/���c�\�D��d�,}��%�QsR��W��^�r?H�i`O�rz��a��ͩ�7K���cC&�o<Ü�]Ղ0���j�{ٯ~�u��5J�����/ia1��EcB�����s Z�^S��yxЕP>�e˫�(r�Q#晓��2��/?������ħŤ�3\���j�I[K��B?��v��r�3OhKX�ZV��`�[���s9�m��;�������#m(�<bS���t֭�ׄ����N�>��y2�0Aٛ��H�z�+p:����ilӨe�y��%��Q4%�L��(���!�29_���,�SO�[�	+�~D�
��o�s�)f+����暧'�[�9i
�e~[���r+ɑ��Q�I�M�XK���C?�4=�!#N^��]��>��a��k�ϳ��d��"�M|z %���)�<O]Z�]}[� l��-d��M����OCG>bm�Wә%k�Q �"z�]�[ �U1�Ma���/�.@�\[w.�7h
ٕ8�nLI���5�/`�����*4Tp��}��_��wMo�N�͎������9U����k�w�*A��LJ�tI��#��#&is+F��nz��V7�UZOg�����~j�989I�}ScG-���~8h��i�:!8���T�aoՔ�0Khqv(�J�-Ȱ�)2����T�}x}��uR�?���D������$���S �T��L����W��GE��"uxi�����H�5�~��ȹ܆��n�(�B��C��zc��2	���~��C�<�=���6a���d��YY��]��(���V:�|H�a�