XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C���c,w�����O��G'��-�`�?!TX�P�&o^�.��L��1�zǽӲ�ɠcB��l&�!����P-���Wm��&�����맡Y�Je��.	e�\�$ �OzWM��Wp	�q�4rU���	�F/5�G5��VŚ�V|Iv�V��O�����O*z6�t��u�����>F̎>H�q
�p�*f���g�z���
T*�<�֩����F#}�#��ج ��-lаlŝz7r�ǭ��.ѣKԁ*儗��M���290w�oB�����9'Ϭ�L��g���2d���N���YN���V��U��q���o>�� ��x�U3�J���k�~�~�4E2�Ole���#�x�2�p&�Г���	��í�W���$�#�����oR��}`?@�.�ఀq�y������ġ ~<��S��H�2��1��
�;�U{�K�3_k`评v�%q?����;��\��3ZI�E���x���u���I�b)���2�U��J\�t�P��e̶��E�% a�r�"����~XMK��+/r".;ҽVg��zG ou�� ������׽�y_e����#Jf��OiW5a��p�ps��!g���#�PP�\�r�z~n��ʰ<Y���_P��{_�ԟ��fb�bo�6�qn��zC�r����.a�E|��8�|��w�<�ZK����/[X�ŧ�Gk��Ц{���p5�IF�麼�a���!Ymt��nXlxVHYEB    1047     4a0���ɏ��%�{V}���Q����"ٖ[zeI���Z�$dE�!�.�A����ɪ���^ԍ�ܵ,��(϶U+���JS֑n�Adl��%]��Pw����1�K���}��ݧ���"k�5A�?�)Oځ3*o�����\9|=��^�7>#j�l�5s���u� OQ͖����l9�s��MP��F����Z� l���<��{��P���P`ƨX�V92��uދ-�cS�Md��.6�VC�1�[�9�o�Y[��kɗ�s�]k�Y͉���"n8FX�Li�F��*�CS�o%^]�f-�#G����&�bW�2[���r����R22�����Í�&*[EM�����=]ϙ�y��l��%�G6L1a�� t���e &s�}#c�+��1`7��4]#\�3mrX�����
��Z��LR+�Ǌ�wلp�m�+R���M��B��u��ke)�U��O�Ew������J���!�d��o�x��%��R��K�Y^p�A}���;���V�t�/fb�3��Y�[3a]C(;��3�Yw�D8�A�t�:uP��GQ]�M�4S*7Ȋ$��N۹���>O�q�0�l���ܜ=,�4#�5�)K�m��L��(4�ǈ�DH�t8�NN�^��z����E�5�6J�TE�b}�O�Rq�%_hv�l�{�G�nߦ��� �����<�L�*��!�O+V`%�|����F���Ü�z9xFtkUT��F ��Ma��No5|ic�J��7����j��cC��a~nBГ��u�,� ��n�^A%B��ef��+���Z+��<:�
���Qd��y����翊���8�d�n�@K.�%�m6����{q��ݟ����YP���mN;{���v �E��D���)8*z�|؛��j����a>�ʀvn�r&�t��?�Ѵ ���o�G����فqu� �TbT&W�X�<�@ �B;����f]g�
�\<�L�z{%*YL���T���W��t��������f}h6����	-)�f�;��תQ��A���N�G�`�l}�^��hT���
E�A���9K�6��⿝~�a�w�'�?�	*D�L����z��

������ Aܟ	٪R�G����Ҷ�׭�q2�;�/�����"ů̇���O�a��o{���(