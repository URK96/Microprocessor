XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� s�� ��n+ ���Q�$v�2/��N��X|�9f1Z>�>�+�c�>g�I�|k�ɳ���;�ϔ����O�h�[Bn6+��4�x�� !h^�DW�1tEa.)բxZ�e����}jQ�^��6�0�Dq-�z�-$"�}���*o%�<�5�/�W�mU���L���Z��(�ʫˉ��Y�DjCy,�`��8���N$_�̕���
��z�VEI%B=Z���?��̙�� ͓W\uBr|�7�J�Ɂ�<P����	�Ois�ϫ����v�|�a�Y`oV��+17�Յ
�{�4����J@=�[�s�k�� |dɳ��#�+zq�Gyo(_�iw������� �V<>�qw���Y>�������+�O�~Ӏ�+H��e|9��@��ﾥ�T�0���d!��(����z�(��kgAZ�7�����N`7)4�7�\y}"[ڹ����F�8�䉈)�oI�\?������x�Zd!�*'�`��+�"��v%�hT�R�ۡfs>J�9�x|���V:(D.tid�co{��d��a�qR���\3D��uj+��2�"�oC>��="ܵNO����mi���o�>��)��TGb;H�	�Sz��'��yjK>*�	80bX ����v�闾YDB�!>���� ��dtD����Ocu/�f#��l�K:�=6��z��vBj`�䂔N^f�Z�~�[���������oE�Y~+�2ǽ����
Ǔ�����岔{XlxVHYEB    3c90     900'7յ��nۯ�`L�J*�Zڛ�����"��b���e0P��Ek�d�K�����?�*5��Tj� EA�D�4T*��.���!�\#�2�����f�0�X	��4$�	�4zŢ*?/t]v��:�6����N ˆј����#�n�<�.fo���"gj���~�,�����;d�F�,C�;�����Kx��d���em�6��^�l���q�{ˆ���Q�,ŠP�r~���r��t$�e1��Ϥ��R�)�i|��O��������ٽ�Y�@2	��d�?�"D(����b�ʰ"3~n�B��&^M.0��׿�<#
H�9(�g��be����D���<�s���:Oj���tc�s�pE��D�J��1,���-k�ha�e)�����T���=�܎EX���t�$;�hRZ�+��~��UzǢ�)�`���A���gД�M���
'^}��.t����#�rH�\��}i< �*���8-1W�<>�<�dy�Y�� �{D�'ǽ�>k�T��O�ŏ*�,E�e*U��b�s��g��'���Q���7�!�`"�R�p'��R�v�_�E)������p�����}��Ƅ�̘���ڲJW���o���J���
 _pq��÷g��L�`}yF����ڬ�ƍ�)��hM��	����Y�v�8�<j����{Kб�w�GUz�/�g�&�0��e�]^<6��yG�J�������ض�i��hZk�MϹ��n�XكaV5ª��0~�G�>x��K���tfҍ#����
]�?�Te��>�l���?E\�*&�)/"^���oE�ĺDc��(�ݕ��۟���-/E��pƫP,I�.8e�}�䶢2��;�ANl�v{�KI򸻊E9ed0{}�C�M�jָ�����L���,k.
:�*�(/�7��1\��h�3{k�{��R)�G��YY7l,Yʄ�ȑP��X�.��+j�C�w�2�6�Q����>y�[���0OQa-������Q%�Q?Bk��oU�3Ag�"L.��`x�P9D��DU�G7i�J�ݴV�U�	��.���B��R4�O�6V)є��3}�tBN�����}�і���	�W�/�A��x$���z���SG���bр��J�o���q�r�~-�m�P�f��Y�+U��4��������ŵ�F�>[�ɵ�"�m.��qn�?��.���d�TXلv#W�P��'v��O����\�Sf$a1��v�l��WX��I�py�%��|��\�D�zo>��m; �k:6Κj8a�R�J����� ��<<2"��N�$k5gz��/��t�>�(T�e�`�}�^��D� Z����ȸ2oJ
F[��6$��{�"IiP[Dh�g=�]��J+�nq
?p�(�aQ-D��'�q�Y �.��S����G�$n6��0�/�--XP4F��R�8�
ͽ)Zz7���U���(�5���4�A�n�Z��7���*�7n� B�ݍ ��Q��YɥB[kP}ro���i��\�<{v%�H{Sʜ=��R�I	"r�����)҉
��CKa���Op;�t�nI9�e#�2_u��7}��d.�������_���h�� ����2��o��
!�~��Y,����K�IH��p%���ʃԾM㴵�3��`-�Qו[[��7X�"]sG� l�``�V܍���h֤�i	-R�d�ƫ-�@���K��m����P�3��y��ޙ���l0Hs�z$f&��4��@ԓA�5y��n��Sp ��;�3�a
cב�H�H���xn��{I:�с ��DZ�~~{gҔ|��rU�[���Q4l�*�y�\*-���6/�:���|K>Ѿޕ�B1��Ŀ%q�&NZ_L�}#'�u�Ϝ)bT_n*I�H˭��������P����wp�3ɱ�����;�>�@˺E:��YP�$�tn��0NH�y�vgqZ#��V����eɻ
�]r��t3����r�������c�F��?�#���puiLk��:ᘩ%��O�B�1�xd���i���t{�G�07��ws���=�s9\E�w�b��ti���"������r�eA��9`R^�����H��ZW{:#�W/�ȱ�ۻ#H�6�����k&��e��敲o]�-"��*}c�Wz�;D\"d�#��K�<���N~N�v��L.Y����i�	<C��e���Ihr}>s]b��×�m���#攄�����]+`�h���
�6 ��;͕G��`a��)