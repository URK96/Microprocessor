XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��p��N��4U��/�n����T*��OS�_���T��e�&�X�n�Z#�S�E5kQO|�ti�e��)����bOB��ke:�˜�y�(����i�;+W�7(���tq��j]����쩁\�B������S�/���)Dm��52�c�i-tn���Rã�7� ���
�d��B��:�$�
"��\(Y�9��W\�4Ǐ��z"�����ܺ�8�H2�m����Y��|�~5G�L]Mz�ϧ�
IoC�S�J5L��d����u��r�#���|\���@	(GPe���l�k�G�p��� ?�z���9'�7�`*�:�H���]Z�l����U���s���+��g�^Z*X!+d�҄"��1TNj,��T޾���ޖ���K/C�#�Njf#�D1���-})W� �mORSh�UZ�0Ԁ�v
+�A秄T��Y�Fd�ȏ<�`ҽy�7v �<�4�R�%5̢�&ݫ�짐l��1(	����-�!��z$J��_6��yz�/j�o3�zl��]�� �e�v� ���R�:�6N����J�?�4��?���'1s��P��v�Ϳ������r�\�&���M�y�wyH�|V�0A����.䰼x��1��6��(���$�Z`7�V�E+�����$��K����1�<���by?\��u���X�3�T���l(!{�F�l��z���������_�>6�ĩ��fa@V���b�������( [%u{D<�'XlxVHYEB    2902     a40]�e�$�DOӎ	�z̜�*���������C>��ᰴN�9{�d|��Q��IQ�N�X��0���,�A����'��O)��D�d���ecc����BY1�F�9y�h6ݞ�a.��7�Z�7���U��d�"499 ?�U�rp{��3��t��T���Zk��1�B26LP���E?Ѫ�դ��F��K�ꥷM�[R4]d����6���Y�DP��Q݈�����U���ĉ��eB��l�=^k�Z���~y������4BOʰ�iPU�j�{-T����H�~�g�ȵ[�����/ҡ:|y��Cp'�f?v�=xԀ���S{�Ƨ���b�%�0���E�>ix�"*۰&��Ӧ�H�Fwk�c��`�����4X����/Z=!9�( ��p�-�*�&d��5䦱��	�=��in�.D�[��,Y��<��`�=����A�����D��nB1b�W+1��u��^����y:ݰ�߇Zn��z+9o�v/�[�D�ri'��Zr#�o�@Ý_"6��s�47�Kg.w�٤�P[ۄ:Y��g�R2�ҶXX9��n�3���ɋ�M��J�Tp�hI�Ү[��:X�3�#e��y�
���!f.$�޴"�㉮L��U���!�2��9���q�H�G�xB�o�>|��3-�;5B�@@��y�n�M�S�N�M�l�;��iq�>Н���q�{��+g�{�!
��^�S��Pŏ]��P=Np��2O�I��9���; E�����(iLҟ���xV#knx�2չ4�q%�!Us4������5��=�YT��ȝ��6�+o#q6��6��D&<�r�|Ő�����gKv��&��V��D�l=,����	���G���y�\�⊘���_������)�<w6��'gkq$瘑��_����Pkb373��/��!�A�Xvώ���Ub�E�WW�[Z��o��=��Y�o�ə24��p^`(�@��&���%�Yl7���o��ĭ����5!�oԎl:�<�T�ʢ���a�-�B�Zw����rѽ�v	F�nh#��2�d�C�<�C>�K��:4�-���(Q�u�=n�k��}ػ9��gza��h���[-fA���3���*�J��~���02�����5�}ĜB`d-W	%�R<�!�f4������*�B��=y[����g�(Qc�K�[��)	��7yՒ$���o��tyZ�{��D�P����g���l����M�Y@'K���Y�F0��!-F!r[����VoU�q����݀�#w��� �9�R�iQ
�
#�x���;o7���%+��>���e�w0�[�_���	���'w�;~�琍��Kp��
�O\�
J�6�y��>��ߧw��}��p�r2��3k5�djn�B)��d%$�����X�N�/ˈ�ٜ����V��>����;��Y{�Ba�;��7�����.��X�������S��U�#��D&�M)�av|��8�g�� F< 
�iq�es��5D����}Vս�����ybA�EMu�F�`!�B�{F���9���!�a��W`OB�Ȼ�x�����n�2�}%A*�)YZHO� qv�%���6���8�KĨ��YW{4y�����ʙ�X�eY�W}.V��&V�s��."��Fk�����Ҫ���4�����/�A����6n��O�D�z�@G��ܳ'����n4�r)R/E�W,<��cD����Մ~�5���C��5y�SE{(�0��������~�2^ݨ��]�l0ٗ&�b��Ox�J!]06d�h�T��.(DdĈ��M���Fgd�K�\#'�e-���$�c\��ܛ��|8Ԯzf�{�.;��I���$�D�p���y�Fbs�vRNLpa\���oS�[��0�7%��lQ��#�.�y^x�w0�`!��Ssn�fa}��7���ϥ��K��瘯E�ټZ�i6��Ë�p����SԴ�4�C����.Sx�R�+�yO���#��W�+�)��ol����S<����J樶h�yuLj��HN��ԭ�o�k2/�AT��)_NF�E̠&�Y�UjN�e�r��~�ݪ�<���������I:����"�I��tT�M�����F�gĒ$�+&ib�*��Cm7��O��� ��g�5m�(� ���ZC^F�  �l����~�;n����>uhC�bw�%i�m*>��Fb/4��'#P[�v�W6���gs#�E'��������}P?��W�F�\K:��ui}9��X�v��̄�$%ȹ�NQ�gP��専g�֩�' *J:l[+��V���/Ԇ����`��%ç9��I����11���3�t�R@��W���}G�Ծ
Y�ۯ^6�j����܌F4/��l߉��=���]&VJ��u�P������XYg$�	V����߾�7,h�S�Cv�Z�����<tGl����?l��ʌ�*k{X�ܳ��@�����9�{Oc�{,��d�Ł�:i@�Լ9��ޔ�XLK�=7�i��8��枡{�8�ӝ I��.�y���KP�W0�͗F�r;!��`�f��g�p�"|:����K�3��L8���D��