XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����8�����ՙ©�W�q�k���i��$�E*q�ݰQ;��=���"M���A���?Kt{�w10� �p��ۤ$>���#��N���W�������
���M�2��Yr@���p��28~h�)��}!%��ﴉ6�p�c-��� �7"�fM��l<�� �^�Zi�j��6�ukW2~��Y).�d�{W%�	T1�r�:cMϐ�UW�+�4Ӄ�`c�k�騫���_�V�E7o���v{����Z_��%A~�H�=�;����뭱�Coƪ��V��ƧJ�*@�3!�w�ѯݶ1����d8����(d���j*-��XXe��*��������Q�
�()uҀb�x�
�Hh]��p�&�������T"�%i`��Z�͊A�$�udbJ�)̍� J�R5��X�������=1gsF,��'�#B�z༦��d�E){�Tf��Hr�Ҳ�d)R����k��Y����9���7���"�Ф���A԰�%��@SL	X"`�T���z-�W�ǺK�g���
�{�ai~�*¨�_%{�R�x=�~Jl��)����c��&�p��7xD�u�3d�ȎE	59P�� #�f��.����I�l5�z��ʌ�1ap@���Un ����RcF�.�$m~��n��w�Z��^�k������	cqb_�yt�hg`a��3��� R$�s��;>.i��?����|��>e�2\���M�N���}��I��E_H_�N��^�<T�	�5�sՒ��2�Pq�G7�����@�#XlxVHYEB    10b5     410���M�.��|�o��k�.��������A���y��C��0)K5����(3&F��I�E�	��Dxa�A369-�$�O��W�y���P<]����sD��H��n%�BD7�SY5��ݖ_�?#��;F�'��]����;�?���h��N��_�4Pa����cu�!ͣ
x97Y�hY1V�	�L��Ҵ�=IT.�D0[� T
KE6�Tk%��m�oK1����0-���"r5��:��+�(K��D_����ԝ )�K�d(��"DJ������Vd���Kl��p5K z�/���*��>r��źp�C6#�'�����4��ɜ�	�ds.b��]�3ܚ���V�5Z���n�F����y��+n5�S�}�e��X	�y�Ϸ��hx�o�����1�SE׌eOtr���c����ɼ���m�U�fC����>�����Q}�8 eҵ���*�!"�w�8m��ki�X�@U�����Kŷ�p�;�e`��]�@G��S�`t���!��Nk��y\L�VjRWy�(P=��)F�Y_����@?�'y� ��7w��y��1�i�X�I�����1y5�5��~@�Ʈ�Z��X��ų.�r>��Yv���8�T&�L��9R�7����fr_pR�.BZ���xh�j����ó�`
��P5 ��gN˓�A�x�N�Q*g���|�N<*��`S"a֘�2������s"h����� �:f���*i�T��7
��<�<��$ZM��KB���O�u������+�%^�����%��ew���Au�.Uu�:���8�̣�BR���:�0��XgL�_�s���R�CN�Hf�@#I"�ޥq/��9�>��"ߕ��@�g�'f��1+Q+#��*�/�V� �k�8�"���6��(�A�$[��pX�'#~v� @$�&2���5����$#�a1H�h��XZ�*����:��pd'�Kp,��S)��8X�~*y���T���C����mBigg��qN����G