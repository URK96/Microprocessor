XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���qTl���.AJ�M�y2؉|ײS���S�BQ*�A6}
�H�L]��x�hm�y�$�:�9��>��w�2 �8�:ʩu34t�+y�&*�|��q��B��_m��$���d}�V��',O��e�T;%����ڌ@�`�\Ƶy�:�:�3*?̖&�_m�?B������rUJ�����n�UNU�~��DT߃�Bz��8D^�H(��kl��5�y=��G+� 'N!�,�d��'M���kj���������ZH�Tj٨*��V� ��ˠU��,�o'|Vp( ?���#f�TP�ȟ�쯒��N�I]9[ň�N��"⫞��)^�,�OqiǏ[�\r4Dׅ��Ku%
���ֳW����oh�׮'�' }HK�/�%�s�J����-�O�����O������׹�޶��.q�W�n䑎�r���Xf�f���4xBd �����H6�%X�׿��]ٱr�*�ϭ�l�LzAX�	KW�9]/��/(�W��|�)i�9�_�5'h�ȋ�����T��r�TX����t���UѲx\yn����{�[���Cw��A���7ָ4�e*C�0���D�g���j.+iQ��Iۄ���9Erb����˗��؈���mLo�jJ�4���nLg�{��۶GǧsXk%)�U*��D���|ύLB�1I�`��ᱶ�*PQ{�)2���"Z�5r�����
,��-(��4H'd*f ��(��g����u�a�=~��5�|?:[���(�\�w�
�m�����&�XlxVHYEB    1041     4a0s��
���\��is�m��� �V�1j��!a���t��Jv�𗤖�R%�2�u�:��\�,��~lz���Y�K��o��u^ilz���>v�� X+�]&�
��Kăm��M7n� X ��!�7��Fba��5���<(^�#��0���|�/b�ƶh�9_,`�:�V���"Ve�	�L�4�1V�s[�BB.?��Nm���|�{<��N!�W�����*�kM���'�1���-tS����2�����Ї���t�K-�R�o�;��-�Ҕ�����.)�N�ĳN�H�,Ǉo��B�>`��"AQbS��r�l��+�2L�����3��什8�9�.ph�Nk��3/���VQ*�h��}@�C`R���+�.#�(��|RQ4�L�a�B��^���[�-ܭ&)�&�.��rE��~��*޻�YJ�g����{f
-_>�b���O��H�F9�̞�Ɏ���| ��r�]����@�.�ޤ����7�C��oH��H�is��3���7�f��3oW\��N��O�vβ5J'�.}�o󞜠���f�-���g��#]n�XR��yZGc2y�2�n������c��'Ƌ���b��k-�;��Օ�C���N��k�:G�ϛ�>t���O�Ľ��F� �PĒc*$���R��ܓ��*��'f�]۵��.�!k@}�.��w��Ce�W�������nbL��9&���լU�m�z8�̻�<�3�#��"����L���)pi]L���|���,�X':Dv�s�E�4��zv�8�qv��,ܸp`�[����pj�b���hW�̙��"G�<��߽�-��G%O}5�6 X���%�4�k\D����p.���2�'��R��ę�+W�%�t�+W(q�49�̟�����.���& 5b(��rY�_,G4v����1hB�x�\v{Y	-�������>ʱ�D�6�5g�G�����U��X��:ߑ ۔|n��Ĝv�ҵ5�1)�Ÿ}��|�V'D��y���v�9�_2�u�p�nH����މI��)Gu�dv�?�t4~�/��F���WH� ��3`e�@Gv�^����=�$|�^����+�b��>��<F,�i�y��	tH���O֜|�V?����Jj��:jx��>���iw