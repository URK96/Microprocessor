XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E"|�+�3�x;�ͨF�!�|j���� ��|����T�ظ�UXू����&ܲ�?�������p�,�NOs��g `�~~��*��q�V��_y*��������\�+ND�vu	�50HA�YP�;���%\��o�?�1�:�AUi���m����Al<b?�x)�� WD��V�)GI�66`�b�$j8����h�Fw(�8����_�y~��@�dN��(`6
�����Mԧ`�Ӷ�a����0�0�u�t3�����+/"%�0�b�F�\I�z��`J�q9\��a� Յ�O��+~�<��P��HU����Jz ��Djp!������jk|�3Li�<���&�������&oE5��)���U-e:���D��ŉH���G_ �a�
���қ@�]̹
p&�而��I��s�dj#>���RM�|�	�o��d#��KՕ#���}GZ]-����J��!��[D�:���2�¯���N��:���������ͮ�9��+/i�-�N,B���:�c�zPv!��t���3�93��Xk�������-�rdg`v�.�Y�M�Z�4hQ���7�i�/����eT�h௵�s��/X������&��]t\`)
l��I��=!N b��.ɓ�A��W!�i/#+<5�.(�����ᡚ������nU��7��H�� �N(��Fcݴ]���>O�ё2�5GX؛��&�YT��)�Zo���6�bY�駪-�Ww`�ʈa�g+�XlxVHYEB    41c2     c40	���є��N��?,Q�;��������&����o� �CN�O#�ֵ/���ț�iE�m�Qd~\���kVV��� ��i�1]2gC�D��q��nTZ6_SIn�2 �n�Ɋ��h�Ǆ��A؍�I�P@l��8�0�n���CF��K��]���L�`����`!{��K5�$���r�p�3�����LP$^ZB�EV�c���oP�9��G��|��Ll!GQIl�/ZفIv�RWT�d�F���h��tK�\��
�#bT�8m�9�jE��Aʀ=�5�¦���^O���󤍺3uf7��6�����C��p�]No����wI��<�˦��2ս4�o�#'.�O��#�5�a����*^E{�gcËH�Ǝ�˄~
�tJ ^h%X���0��k�����#=z��:��;,���AJk����a:a��H������C�_����>[*#U�䨐�lG*a/�2�> �<cj��x�b3�O �]Λ��A�W��8�����Ik9��&��{���*86��Z�-E�^�#'W�6h��ci�Y8uҟ����u�>3A8]	�:a��ܱ��B�F�QFK:L�o��\��-E�gj�i��h{���	 �^��r��-k�n䤝�P�_��5�;}|�9��{�M-��v����v_w�����п�"��z�F��gI�@�z\S�oԘ֗PMp��ɗ�-���9��ݭ;��h1�S~@(g8�*lO�t}앶ⴅ�Q����32�nZ
����w���-HprV���_������ ��מ�M��q�7&����d�l��U�O��շ=��6�!17|����r�	��g�
Uُ���U��I_Ğ��:�o�3����\u�!���n��O��KBz���}��,,\c.���<���Z�����ԟ�b`�3��׬��g�u�N\�{��oW޾{v<g�?����_0��9�d�5�Ub�F��a���v-fT�͉�V���״س����b&��I\�����gp��K�0=4'\�i�ytwBvF�>4Le��B0��0e,dKm$К��S���N�Q��Fe	���(����{�)]M�� ��Uo �࠽���:�oS1�޲��>Eq�
��v�n��=��zq��a1�7���C
u):� ?�I�,��m�b2Q�[�����2�俉�%� ��Y4De�`~�jk��z��,j����h�k���w�Vr��/`U�5D��g�(㻢�<dGk�An�O6`�9h�t���I��=!1S1m�?;���;�C�a���H� ��,��w���."*YSV��dgx~��$��&$���c1ɫ�	J��;���W�{��T��j>��A��?�w@؎jJ�
$�^�C.��޷ l#�3F_�lQ�� KS��
�h��;��q��[ُt"���VT׽;��ུs�w���>�`c��5���n�.9NJ�m�t���-˄�k�\���h��?_���v�Y� �8_�Io+��`	����࿄�^céY�rpW�i�F��!,z�Z��-�o�ca��T~e��@h�l�T$����P�����н�{�{.aq�[pDR3
<S8��#����-����!�_��x�Cy���1��R�����K��	;�[�hZ�q��}8�_h!h Mz��Ġl��EU��Wv�Z��N݃�Wç(�cS�Qr�5�T����o90����e�I�n
�˝�J�x�X�i�V�LCu�l#ݭӫ�ʏso� c��Q��%�+�Pc��/ܿ@ b-��G��r=�K�x�Yʳ̵V�u��j�h�O�?��bO`9M�rX3̇~6�{D�ѽ/I�0�_@|���IU�TVsIN��d�j͹�/��+��ѱ��h���q�z/u�O���[q��\�g1�c`�Y�j;�j�o�DJZ*�V�Tm'Z�r�˖"��[��kܫ+Xf;#M�8M�`ܒmV}��D[���/'-�e 2�/��utn�e��Sl=�J���س��Q�>��.����ϵ� O�C�GC#�0��1�V�#���`+t,3�x�@]3�傂�}����_!��$	n�-�i�#?|��	��)�P�x�J�Tp/'����?2Q�zj�s�K!S$�"Ք�X�-���ޠǩd�O.��f��!+�c�@&��XB������i+ǔ�)��ǿ�1Q�<e��qy�WZ�G8�=|]�L� ����X�^pES����3ܢ���k��w���.��O�Z#����{���&��:�F���W��������v��ӴԘ ��[|:޾�X
$E$[d�~�V�-�_�e��d����3�[�޴-U�S6�e�*+���q��#���V1�����#�3��=e(��M+�����j+��b��,N��z_���ò���jc9�{W�u^����E#��7�lN��6@�����W�3ZQ\8�*�[?���=GV`��Y�Q����Ab����)�ߒ�@A_h��Z�DbX��s�\�(c+C��T+;A��!9�[����x	_�VV20� �1�0�wm�l4Wktgpw��=PWǏ�w#�Cf]k�L$��GE8ح��߂�E
��{Dt��-ɽ�-m��o��RTe���,�jT{�s�Q�( CمD�A�4=ŋ7�g�`V��;�������[�0+nM�Ӭ�\R(��Yj�,���� ��=&��^��������s�}�E����*�řբ�9����D�0J�����N9�M��4�q�t��_�L*�s�?)F`���3g�R?�I�?�����j�����␒�h�N#��^-t�!O��������%��b�`pzI����y0�O�l^2��1M�BމffsT�S���EjT<�F���j^�hx�9��8�-����%�G�y�'w��`�TV�5�^C�,h@KȔaoDOb�騪�4S\��~S=���`&��(#��e��eb�+�x'�\b�����3l�uc�X9h��������h�{���\�N�����w�
ݠ?�}��p	���Bi�-��J���0��Ш�j#?5�Z|�ws'����Z���H61ϰ�o���f��rU�Yb�k��#�O\�ֺ�p���edr�mC