XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����@& �oԋ��t}H�������D�����V��}8A���=x��?/�clVX���C�b�r�q͕P��'-����:c�#.��:��iD)<G��Wqׇ��O�V����	.FQ�����\���͖��C؉���]Q%_��ŗh�N��4`h���R���
�.V�!=��**�C5�����n.ؕ��%}f �0�q	�����"�@�驃v;Pm'!(B�q2r[��	zCڧG�ʻ2L�ְbj�|1`	�)��T�=}0f��9��$n�Zp~!��8J(?��g�mU�	9F�U�C q4I86_�<�b���`����/`���G�7�(٨[L�A#ѻm3KJ�fQ�P�8.�X��1S^4�E��F>�D��035�ـ2��	'�����3���^��i0? ��n��C͞YZ�-ԫ���� ������D����u�K�{�b����݊���.�x�מ�1�ԝ��@��`Hi�k��M&#���z*Ec!��)�ze���]]����}���Fu�թP������#�(��?���{$=�.�zaQ���O���~uR^-�;�WDr[����g?*�������1�gD(�jWg�E�eh@���J鬠�'F�)�E<!�ŹWد����д0|�"�������^�s|�t���{��߫Q�
?�Me�(f�el����V���B�5�8���|�R���C�a��H�����d��
䵛C ?��O���a�q3�r��["�"$��XlxVHYEB    1621     410��;v�!L'��hh������ �t� BE�����	�y�o��0sc��2NBzH�x=N�9��ci����^@��-����k� �Tm(0��v��M8��e��I�� e)-�h5���,d���'@Y��/H�*�EI�ThW��+�*a]���@��7$Z�`-��d���� ].
%����Y�_$�O ����$��1gt0T���P�1�}v�;
�΄)3Uj������� 4f�7��i�
�%�g�XJ�!9I]6�S���# \�,w"fb��ls!��P�ϧMʟ�6�nsj�~�F��B����$A �/�HG'��c��]��
��&��9���:y��v����5�͙6r�F���<w������>����+���J�oH�0o6�\l�h<;�b�+b���%1�����*#�)�F���w���S�Q�}i�i��u]l�
���XR��ޮGd֓���'&_Y�/�s��9��+�#�m�Lz���y���C�d+H�%�6s�TN��w��]����?/3"��Y^���Ʊ`�!z/c��SV���x�G6�7��"��g����`�2�h<�EN��ߘf����u�����!f]�;`lnF��H3Q[[,c�j�k0���?�U.E0B�0�I{)��&[��7����w���JE�������U$_h6������%N�Pe>�	���H�X�L�w_�ms1�e��:#��~O��}�/al_�^�a�A�!�uquڕM�#�\��,��R6��+�X"\{�/͗	A�ML2��o���c���J�Rޡ�Ȧ������|�0��:k�aU�(U�Q�7�g/Ȝ4R��q��f|���"��v.C�O��9�P����L3W�X��~�ɒ��bう��H��,��@���d�a��j�;���b�p�_��%o(1\Oؼ���8��pLI+����?[ztB��Mf�`4�q:W�UY2���ȅ������ǎ��K̂�n�\�Zs)O|��KQ=7��	V{�D�:���ej�Y�"��lT