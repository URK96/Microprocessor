XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���p�'9�gl*�&Ā��j�#�#/{�k�܉�1�O�2��!�ޗ-��O9K�3�K�o��Ǜ�?ǘ��l1�T.�#%W`�$��s`6qT����s��t��L{��8����L�L���8��لA�Q']��1"E�DxWM��d'/�9��=�Y�țM�I�r����;�5���|�j�a�$9�/-�������〲vC���
�F��8�R���;�7���Y�v�w��;~�%�&���J킺ǔ�>͂���fCrQ�%����fI�]k����\#�9K#@cmt_�L��^��N�rBtF���pZW�P���,�[�����e ���b�U�� H"G'���0�+V�BkI�9!S�;_��~YY�T��6���j��_n�l���k�v�Hu�A�U�Eq�5A�;e!�2���75*޲�O "k���f�o�I5���
�y����,�C�(;L�0��(ѿ��nq�f��/
�,���[��@{u����pT��y�-!	ƣ+*>z���6�5�w��i�vrC���U=�����q� �m�$�c���5��,dM����)�P>�f�4D7UyL�C~��$l�����˭>�@�$5�iq�O����`4|j�ޏ���`dj��R�U�XupY��劣YM"�u��e��b�}��Ñ�����}�C4��Wf�wԉ-�!訐Q�۹��↍xaE/P���
�"�j��U$Lk^�'��W0t�o�
Rrf�[�8A՚T�^/�N�cB�XlxVHYEB    1d53     7b0x��V�7��b-��X)N3�+X��*�{�Ĺ��R�k#��&���FȄ���3���Tk��f�vh}��~Ha~��L��1/="4����-�$�t�'+J.��z��W�O������>�>�C�*�ltk�?X�J�IbU�T�g��:%(�w��8��~%���Mi�_�]��ș�9|��<H:~R_��1y�5?<�$� �[r�a���(��K5�;��[?岅�=��A��X��5�w��N��<i���C"���nߞ�t����^8cb�c�L��_>�M��Oo�����k�gE��&_�^��v�	~�՜�<��[�ۢ@�p��~
��o���)�|�x-k��T��Mv�$k���$�������TxB��\�ϗu��_h�q=�:À��96f�/f)0c�?���\�y����/p�z��O��Wќ?��S_���'���J�r�����_/H'����Lh����w�#�;�����Q�����y�q�wS�HğE�n�D˜���#�H�X1�������B�&��(����yxwDϵ���9�{�y!��%ə�ͥӻ�,4��t1:�Ğ��b3c`���܄����}���$<E�'qAy��'4-S����h)ۊ���j���o��hYu��g�E0�%�n4�st���@��f1�]7�x���F��0�T^��3���G�SV�?J��h��}XT�;���a�������Z�w�`����އ5�&�ӃlVv=Ӱ G�w��
{���x޻�L	d���GH�z���-��h�k%�DW%O��s�v����	�g�MR���[��0[5-"�6�Q=Dz5!��Bj4����z��=���Ȯ͹���Ѩ@�������Ƙ��;�� g�R�F`��e����3��W,\����JI�v�W��Ew��MҖx��E�/�7l���yz�k,��H�_0W�UĔR�t� 	����u�z�F"VL�f��ɝ�_߶(7N� �5Kv�ұ��{�Ь�vPxA��D��eO:�l��|�o�AF��yF�܅���Z�Kĵ(�ǫ�ʅ��m}�qN�����;徻����k��v��Է�_[��%J+�4(�Ot�	�6||��aDt%�"A�*}�M )" oy�kc����W�E6k&�����v�G`����nbұ���4���Ou��B>$s�m��Vx�|�[�N=Ň��~�C�KY���Om<|���NQ�uc�Qdޜ��Qɖ�_==�o,���V&VI�B$�@>,^q`�<��zo����O��WuV�+f�2z��nF�n�ʖ"c�X��3�/ ��)
+Z�9�r�-��p�z�j|����ar���Z��{thG�ҴD4�
�{5A{1�>�Uz H�kKH?�S�-���2�(�Y+���Q�F�F֚�^h_���3konQn�l*m�p��0ot[=t��)h_���aE�HҺ0��j�JV�b��s|�D8C��y����笒��(���{������^�I]m�ǸDϋ�!�%�,�)O.�P==\�ΰU������қ��^��8C4���hh�D�a]�c��dg�B����̗��Q��.X=q,���0m����o����r���<h��qTT$�&���rN�v�՜�-��)����{~Ē+��6���R%r�u(�I��6��j&��Nk�g����f"���ڜV]u^�H�}|���$�v��;kW���k9��# LqD+������=�&�r�Vf�N<>DV�[�.0@6}k7��\�.�'�����A,��PI��n�0]ߪ����9�ll����*�G0|0�������;Ť{<W�z�� A�W�3�F_�.�����o�}����B�
� s���r����>�㯲��l��� G�ԧz�L7-���8����Om�%I�y��R��tSׇ������