XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���8�563�D���<ayn>��r)c�����{Rm��kB[�u�>�@@_eм.�6����Id��$��4|��7�qQU>�>���A�}����`܅����&ha?�j�,UFh���:�c�O�귭C��1�@̛/Fbo�Hб+�9�?J͐�E+�[Iv����QP�4F K��<_^V���)z^a���pj�	�+?��/&2��Y����*Eܘl��t������c8��Qx3/`�M��w���.���zK-�@��e$
�;�h��H��q�������?��7_`������
�oK�j����&æ�F,��_2 �2�9��*��>X����S�߰�}�kq#ڿR�]���'��"���)'.H������%�a	�`�,}ϕo!j�&#b � �p�y`��AbQN��a~�h���,���K>�u�MI��a��n��CIh�\�����K��]tΆѻV�������Y�@--o���Q��A�i���Ë��!�L�zX��7� $�Z�V{h�M�H$�u��A�j'B^F�M(2�S�a�K��*�wns��1p��}9l�T'�]%��6�R���}cn��jrI��Oq/�j 	b�/r�&n
o*� 8-G /��i7����eI^ϟ�Ӱ��F����²�kb � >[��t@֮�o�d�F���?"� �?p��@��Ò�0�:r���-*���Buo���P��}�EoWٿ���h�w�V�⋸V��ތ��XlxVHYEB    6fd8     c30;�(m�R>����w6�6!$XfL���_��T����b9m�@JCQI֎�Mv:\����~`PP���_��y᱌*�~�	��LF�q�?��|!��K��Јx��~R�iML7�`�:�q���!���N�sw������	w����r�}�4�ޞ�Kke��ã	���]Q�X.k5�`�����e��i3�ڴ8�QA�A�[�jζ!#�]���#��g�
>H�ygJ�y�,b��y���c����k���A���侞u��ѕ���vX�x<��2��nO:�jT-�L�_�v	�.u��6�#�ޖ�O�N�-�ٰ`f[@�5���nTCFn����t�#��J?X\�6N�(���Ub�F��(�P����+�3����I��������k.�rb�����aQ�u�YYR��H=}$Ř�F�w����ym�p�G��A�'�G;��ɱ��Aj;l���M�	���u#���[^^�D ��������O����IlEf"¿���}z	Y�������X-N�T��,*k�ؠf���-�;�������5����ƒ�g���6)t]�g�����ɔn��F�)�p���cs����,�q~!^���~!Lfy*��kKF���*�����d�3W1x�giN���"Վ��쥘��H}�.7�6�"���q�&z�e�0��f�
��,wZY%����<(S�r;>�U��۫J�wq������)���ɯ�E�೘"`����h����P�0�c䠠�_.+���j��e�NdM��4[:�|�����v�~b��욺'�v.>�{�G5�h�Ie���=nw�\Ʀ{E؁?~�è<���T�|.�4[�ą1<�U�d�^��E]��쟖�c�"�"�\Wc� ���?���Z���̖�r1��V�l0So�Ԅ!i7j+�������z	|H��-�[��A,L&�B�E���H�|�aP���at���#Ѹ{H;c=
�*}CL��K9���Q�'�A���i�Z QI�F�� tv�� 7E�p��tt��,p��Uu��'����"�wZa����q/d�E�)'%aT��'�J�V>�A�=i��q�^3c�[�g�Î�=�=����0�+�,Z��H�3[����V���[V�ON����ŽH�ߗ��N�/DA�w7��m�%w� U��P�0Ľ���Z�����sPϬ6|+b?Rc;��ać/��CX��(}M��Z�U��v���|p��]01��m��E�ߘ���']���x����������^�JY0��5
�C"��< ����ӂ�}LVD��Ǭ��+sF��hJ�7�w��̓�,�:|X� �W����I�bʦ�j�0�V|�!i�z<۳�����Hߥe
�����T��i:��,#�S�ۭ��8�Ģ�����#��<�X�^�[�n�_q&�sj�Q�9�U�$��=|6����#:��	?��7���i8��u����P�T��QdYs�Tj�n=�4�3��$#'�)�\9Y͢����>�lJ���I��w%�N�����O�t��/8��|�C��.��n3X�}"B�I-AQMv��폊�e�y�0��j�=u�����9C��
���@�).z]�;5~�}�WѼ{�b�d#�[�{�'�Z��Ӂ`��\!1�S��ӗ6զ�`>�U_wqԝ��r�=d1��� Ga+���VY�$M���$o�É�<��{O���BKw�`ke�À	�ϥ����d��������f!D�:�/E
D#�nKua�SX���P�V��̘d�(��L�K?(�Z{�L���hc=�WK�¨��t�#C�mJ�F!�Q={QF�i����<σ\}zD�?�m�W9��-���D��B���
��m�gg�-�|/�,��~@�*S����G�[<��;��O0{.��5WQ=3������V���\�I���x�S�yl�V�9=$h--&W(���u<�q���J�.��D@��(�!���U{}AAW��H=�M�u]/W'<E��F&��bdNܚ<[H=0����\���F�A��^�@(\�4@����������S��8ܾ�DF d��^�k?K|X��gķH{��Bi�M�Yn�HӔ^�����H���)�2���7NUx��D*���0�O���E��U�N�j_��.�5Џ<_���T�F��B0Iα�z�%b:P���D�  ��x{:���B���G�VB����.FnW�("�"s?���t�`}��f^I��Jş5�>�Ԏ����k�>��/dJ+���H�XSI��:�$^	�I�qb�n�t�6�U��A(���tSGBK��G
�C��<����qUd�#�����a��y���b�[%���H�ł�銋�Ydu�u�HH�Y�DD8kH��3���xu���V4��٫���5YI�6XUFNa����|��J�<2Hlo�G�Pp[?>ۮ�-���iW?8�Ύ=E/U���p�	a%ڹ$�Y_�Xz�GZ�
J�o�����������nT���{0tJ�rD��uhb��Ǡ�1X�P%E�m{���g��JQ]����T$j8k.��΁�W���I�K��2sm*Z�̹ط� �ȯ������@Ce��RQ�-�2_ǁ3��P� R�X��-��'V�2p]9}@�_:D;�2o��vC򻹉���"g |�I��6��my~eh��w�2�܄;ZA��	1>[�
�v��@�KLځ��@*��Ks��Vm>�Ӌ����[=��:P��e�`�L�c����dA^9�;�C��Bb���랓�<�M��&�]��r�����~)���6�.ν�ގ=���r��L��|������=SV�������������*����{~R�%�{�5鴸��g��6:�>�����,�*��Q-�m@�������!���5hDF�8��
O��a��0�|-?j�_ÞWD=��[�`e��TeC͂�����52��c���3�K��K���ǟ���J��+�>BH��_[-̝r^�p9�y�*�O��M	��Zk8'�
wؐ��