`timescale 1ns / 1ps

module ALU(
	input [7:0] OperandA,
	input [7:0] OperandB,
	input [2:0] Instruction,
	output reg [7:0] Result
    );


endmodule
