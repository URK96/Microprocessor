XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��dDH,�)�q�<�1�((-�1IٹwHY�3<9,
�)�BylXc����Ke�F�Q�!�7o�F�*y�lr�~�U�e���N�~���{���UC ; 7��G�r1X҃Y�.��h�hxw�]�UK�ٜH�m��LQ}�5�0��i�T�p����T�)`�;�x�BH��A21��*j�$I���t$���$Ew�G��j`���H�y����B]��6ٝ4���f���C.�����Ɂ�9��Cy�߬M$�u�M�fh���\������Or��L�=#F���5}���l"�����5�<=�.L�m�{&jC\fݼ�	���E(��U���&v+�̬"��@-� �H�N�l�p c@^��a���1��507�a7;w٥�qlܵ&Q��q��y�9��*'���
1��F\3~%tpV��\Li�8�Vd�1*/#�7r&�[���Z��-Q���������㇔ǁ�\
��O��`t�)���Ж8�ؘ�/�ۚ�!�[~�%F�ueNN����R��pSݼkNhڴ�I2AKR��.�g���S6�m�����=dY��	��
�5=K���WxE��L���
�@�E��v���M��RE,�=[eXJ�O���|���7�	��#7��������Y��q
a�̾��	�uѰ�,�b�z�>+wpwM���Y�=�ˑ�Nf���o�ʲn9n��E�%���>4* �$�W���m�$v��v.veJ'���X�}c4�XlxVHYEB     a7c     440xfݿ��	
L��#�#�+w�����k�a�^�����f� -�Ok�H)h#��|�Dɘ�=�)�������y�r^��$ؐ�S�d���[��f
O����C�
	��9�4����7a�R�$Sc���p�xUC2���G ��R,��}Sn��_4t�[����qg�$�2%R+��j���þ>T"1�JK����t�v ��n�H���n 6�a�A��3eg{[�c��hO����n3����e�Σ'�*�È�!��(�{�x]Q�� �h�s�O	��C�
��v&���h��K�Dg,V�����W�<�J�B�x���&���w}~�T=p�5��uR��7V"�wn�Ӄ�[AH���ɚ�,U2��;���'<�k�Z�l���-'�a��kS0X��.ʚ�Ϛ�3���N�Ԡ���U����H�i�T�����!���=ß��ABu��a�U��f�6ODK;�)�)����)N�p�*<��+a~�w�hS�_K�����6U�s�T�_�ͻL�
�2����Q8j�ʅ�m���b�R�Aҟ
�`�C�-c1��}�ZQ�����c�j6I���W� =�g���n�dQ��u1R��A���.��v6k?��?CTS�@�\�f�ϧ�}�@��4j�3f�jt7؏�+uv�a?�_u�aLܤaGC\�s���J�+�qyd�-����%ˈ��g��Ax���u&��w3�~�Mdg�PK�"�Rڪ�ׄq��Ǖ���&��&��c�S0�AD"��#�h.��J����M�"{p����ю��Zr#�����.ۥ2!i~���	�J)��S���m��Ui���9T!�ށ�g�eQ��<�W��f���2#�4Ș��C?G�*,�:~��m�=v7..oH$r�HY�ͬ����9�~��Y�"+��8?}�s��#��k�s�lu�"Yy�o\z���gL�D��_X~�5+Fh�Beb>țE Cn��$Ǎ��&a��n�4�4w|���#[�k"�|���H��h3��m�]��N�1�ҋ���%O��P�����p֧w�q���.(?���ᡈ�