XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���i��M��ظ���k���$��;}_�L���:?�z���j�8e�ʯa��zwĔ��J�����^a�1����|��]���(�-�4\i�v���O�'�:(�fS����Е2t}$���3���Ӟ>洄�-��0߫��/����F9�k:�+��i4��k�������9F�X�zșDݽ�;c�t\&���8�9jV\�6$[g���K�G���+{������3�u]�� �4�~G��G?ʖ���+�QI:�4�����䉴��\��C��� ���ۊ��~�,�vOk��'��:���e
�h�x@��K�4Re�2����"i��]����!�)CRQ��M��Q��߸+p�J�����y��#&Q�M&
�?,u��œ����$�C'�}Jů��*��	C��0P���[�3`�Mݴ���Dv��d�-ަ<�b+� 1&w�I/+H�"�J���Յ�.�Z��:[=efK��a��<�&�{�܁�Qa�W��^$�J�%�O9���B�*�6I�Y�^n�����H�k�zK5 $���(��^����\v|� ħ�v�	���EQ�K�������U[��*���R_@&}��l�s�+ �;Dl�^EK�����p�5x> ^[~��ݟ�'�����;��G��UJ��ֶ_���6 �]�s���D�܌������<�;�2�?.�z�ӌڠ[�����H��cw��@���4E��L� ���88��HlY��,P�@٦��u!����z L����XlxVHYEB    1577     5a0�/��@5?т\�U��k��E��B.�X_���X9d¯*���.�ۜ����OjY�[���8O�$�1"H�0]��&Q�ڣ)��sN[�|������^�F�uS���|G/�@dS�q�^���n>�3Xb#�#�&��GE�������lJ=�IU+��h�-\���w��U�Ư�C��s���qRV�BN���U Ɖw����&L�����H{Ѻ��]���.�G�b�`X�;��O{�V��
��f6�($�r���x\�n.,5�7�$�&
�1yЉ�1�,��ʁ��@q�jhx�����V�
��N����$�-��=wY���Н_�q�̴��W��gJ�EpLV�XQ/���{i���l�+�6�Q|�+�L��fO�$�yp��+z�A��G�m�@��-EvY�G+P�g����~�d�r�Y��/@L;]&n5!K��C)�!���k� ����9bq�n���YU0U�1�Y�(�&˾���e<'*`Vݭ3Y��w�@��Q<K�y��N���е��V���Ӧ���`7�K�/�520�0^|�C�om@��I��0���zFH��<|X{��"�FS�o�IZ�Ÿ�|��8�����-���K�0�
�籇2�zGK�Vȶ�ybɛ+��P�tg"��O�=@�9�Ƃ��#���lY>��|�1�����?R$"���Bq��|=z.r���X6���$�bo�b(�X*�L�ޣ�4�׻�����f:K�;3؄A��M� ����;�����T�tT(�sO��V����K��~J;m���<��������b��q�@���f��'c��Y��H����Sn�*���!��}�Ȅ_�(y+�G�-[���3:�uZ��nJ��b��F�?HWw�'�m�2wQ|@�����?��'�
����n�߀���=�n�7 :�<1	�j���R����uO��7��qO��~N�A�ȯ��4�Dc�3�6	E��S��������4��.ŴQ�ן���ՆY���/l\���,���	4]�EC.NW��1���@f�~��X�k�~�q�x&��;�oJZ�K�$��M94 �^��F~�#o�{�O#��><.Y+�z�����1z̏��j���U���N� X��p����ОW�W	(�ľZo����=խ$4a���q^|b!���JWy�\��Xy@�j�9�=o��)VJ�Z/(@k�b�)V�[0����۬)� 
ҙp��z�3���&�+H���ț$ZǸ=�V �o���(��mx<�^�g��y
�`���W�~3wroqkEN�s��>^ű�D4qcէ.��|��/c��yh�D����T���pº	9v��6I��$Z�B��8DU����N�.�ܢ�=j��� S~ 
a��e�.鴬��&�7<����#/i