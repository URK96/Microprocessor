`timescale 1ns / 1ps

module Control(
	input CLK_In,
	input [3:0] User_Input0,
	input [3:0] User_Input1,
	output reg [15:0] Instruction,
	output reg [3:0] State
    );


endmodule
