XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��jʐ@t@�):��p
��C���M.J�����U�"ӝ�PX9�V��!i�j/Q�hq�KBY3qQ�jLhF�q�
���?��|u� u8���0E:&$�����O����R��f�����s�E2L���w(��i�b��|�@����''V�rExLq��w����[^����R>7�DT(��o�ԴC���{u����(���S�@��) �!t��͆ȍ��x��#�x�qGx��M�.�|h�=PJo���Wh���g��tR��l��s$rF���l*��C��C����#3���O-�ç��^�~qF'��8�(7`j�h�g-B*D�X�NS��&�78_�5�B�##zRE6���MK�_����J���y�J���BO��=��Ү@���c�j70��ʗ	���Y��[ʬ�¡a��<0�^�&�x����@1���sid���`� ?�uz��TG*���͍VF�M7z�Vz�XD�ak���wrH�c�3٪!F%Q�X�t�"��"��.@�6����b|%0�i{�r~@�Fξ����4���7$PP4� ��=���7���w?{�����Ks���&j�k���	��L��;� ���M���� .0�9��h��I�ſ4�쓾�#T�1d�Zg���;�� ��ψ �j%��˯;f���Y/~7z�=�S��ƷIy6�E����Q��"ˀop�{�6��N�U��ڐ��A�k��TҮ�W8s������ڠ6���T��RXlxVHYEB    a6c0    1b00N��ݯ�V����*��2�9W��;�P���.�{5��%+K��#E�1������R�0C('�?�GӔ͹��C�	�[SPy�nD�C��4�>�<|�~h6}����#iH.~�vG�5xC�U"	A�@��ktGP��Ze�̫�0�fo!>�ڄ��s�h��se;���׌�Od%q��Deg�
����6��Q�Pįư�;�h���Ժ*����w�U�|�Ȼ�{�G¤���h��Ce���G�L��?'Ԃ��J�`R�8ݹW$��]�IR���2MYl{�
��"���D=Am~srm�E�.y}�H~�=�N�Ok�WG��M�xQ������iS.n+����WzF�7����"/���鑗Q����pe�H�:U�`�ΛI�3�m��Ә6T�/�X�dc�B B���`�W	�����2��7��wb�=3�G��?�o�:�kT��t��"�NyPB�פ��YWcv��As�C�x^��%�6���gqZ�`���g����}�>z��ʞ��P���6#V�#>���%��-U3�,���(�����nH Z5������F|�q:��	�`T�Q�N��&R��>LiV6z��n����/r��9���1�Ƃ��u�,l�ȣp,6�(2 ��'��e��h�t�=��PR�2��zX)
d^�/�����<�s�-m��V�㺻mPM��Qі2�%���_ ����h�1�X�T�eKȵ��-���7�J�h�4�˧غ;#�> MvW������-S\����Ec^&:����' ��cP#�&�.�;��|���_�y*>�����؄K,���r�^�m�z{06S�m]�5��u�q������-���2{���5��6�!;b=���dE[��b�b.g,墸�(���e�^[�;x�����G��^����{�/���Q��2�컧b���ff�QQY;��S��'�<�,�t���UU�m�[��S�EU%�fW����U���F�����jR)�����d���cJ�{�l!�#F�����>*u�m<��v������l���S��8���+C�	�۳��u�	b�����u��:��x�^�Ŭ+v�+�śⵌ��O��A��ft	�\��2�A��?�|��/ :C���v�R��5]b�%��ڧ+B�s�X�yqy�?�>t�y���qn��9@B.�!ىf�
�[���4F��,�ed�B�śW�"َ�'D�S��A�����^[Җ}�2B��(P��cQ.���9 J���W]F�����H�I;���	
����\9+��jah�@�M�~b"��2;���^$T`0\;1�TzL�(<�1���}�D��7�c�3L���q�	L\�Z0:w���Җ�9z�-�xptz�9~^�Pқq�w����~2�6�[k[���sz?C{H!_|4�̹�D��i^�ER8�ê��bp*�~ʙF�&@=�!s�����M�2��%���9�,�%�����v�|PVL��L)����A��6k.�]�<}-T��+��̑#?k���]���bc�5�x17�P�_K���w./�F���x�3Y����:��q�lS�%���{O	�����7�wiE"-���q�z �|zQ�˵*v�KaRu�{9�y�Y$��r��8PeAλ��E0���}���pI���OŮ�O7��H1���+S�ҵ�t���Y<��61�*���.N<]��{�҈)7�q�����s҇%��'��%�;˦�Ձ#謁�(�!ޞ!����DgcK}H�㫻��͍���{�Yc�r��d���(%���ܤ�D�_%z�X�=�p�o��/���=��DQȚ�=��^����3C���2�M�J����Z�z7��p����;�O����V��Gz?�5�D`{6<w�%���u34p�t=�lN5��z��P9�6�	z���!y�9�˹��GV|%�K�/RВ����%��ga �:�6���y�{��%I,�φ��<i˜��'#,��ޒi'��^����s�Q�E���y�Z= ��|�H}����C�Kv����\�s	1��Ͱ�=hQ�6�b"�(�ƪ�NZNj^��;8����*�9$5��y�c�6h�7���Q<Ep�B����b�)9󏎔\�ɶŢ�ͳ�d�����\�=wo$�)n��M=�:r"�[�Ax���KǇ>�KX�/�����ud�r��d+b#�Դ,�Y�"��q*�udXd�E��(=�ރݣRF1�+��'��Bt�)w1�2�� 	�@?�R�ٚn�=ˑ���:�<ƈ��S��-����a�`Gz>d�z�8���Z�	Ȃ�C��V�EԲB̛�?���^|�c�eU�Pt�2d�
�*%牱�?��CG��J]�_�q�)�1��Є�l�q�>H	M��i7�C}���0��0�y�[�D��i�����~2\����oI�:�F5�K�+lN5#�涢��_:n{˽��4
5�Z�t��Go�.����g�虽�.���6�D�T��(x�̅3��<��\b���%�o3
�ge�)�sZg�s������ur�ڂ�nB�]2��D��q�D=�$\T}˝l��Y��]���h\7��6u���iH`��Y�ua\��U����Q��˱;����y��߁yu�e�y�}�z6ם�����w����G����/;^[��FPZ�7r�
����v�ڱ:�z�����o��%`�g��Lq&1̾����s��*�I^;�u�z��A,h�3��{Ҩ���H��A�o��b����j[��.`Z��.��N�9K�յ��xo���[���1u���s~M2�7"Fj�Lqy�|���(P)2�fȚ:�=Ҕ����F���8�� ��0�{���
��CW�~J,j�{R|4d�R�����Y�3��gr]S.�O*M�+��AE�c{��F��@�uND�W�JWf�v�vW�k��30-n^_�~�/��#V��[��z�z�,8g�6�u�������I</�j��+h���'AQ���1�es&���#�㉶�k,��6�
5��h^5��A��NL�W�A��� x���}��T'%1�/����Z>���hq�y"w#F1n/� ݴ+�8J��[�;}W�o[�g�B�G�h�4��hB*�t�6W
�Pd�n�ĩ�҇*���l%�Z���i�%����w���	�E�t����3�O�V�&��k��fw4�*����U�>�\<���#���KS�f������E�b=�iXtJ���.�گ|�"�h����������!�0���ر\^�?�_���*J vSv�[eK!e���@�+$"���kF�������UG��9�K�MH��Kc.��K�U,�l�����qȃ�F�w�G2�䂛=���7z`y��}��K��5D��Ӧo~U�&xaˍ�o��f�Z���Ȑ�[x`��]����k�y �<��@1U1u�L�C��],k¼��JC�ŀ%r.��y�6;�7�%���v')���F`2�sV#�ţ�5����`]zYI>ؾ���~���ؘ�̈́�����V�^�o[��p�pl��j�~@�5�i	e-�\��v�^uoK���K�h������j��A�7�a�1	{X��v�R݅���9��׍`k�p��yxEWT����2ލ&�a�� @�E'�Q��{}�2Pׁ�fʋ��nL]��	�}�z�T�H�|�Gjs� V��UU���NeV3�	G�g���~jݏς�X�@�ݥ���I5�a9
�V6S����}�J�G#�3u�3,E��,�X��;�Eo=�k�~J����x��-����mp�ٿ��}6��v�^c��&^�H`z$��s���"MA�$�[���e�K�)�����.�Ӣ�k������z� (Q�������q�Ȧ�$r���CEP�0�͞S���]GvW.���s ز�2�xC�<^���/����K�n�<����� A ��o)O_IxI���ڬ�V_S�g�9�tߍ譮0�{�o���{���zA(�J�Įugᯤa�[����\.3m&�E`��2 @��4�8���o<- %�rٝKo�&7�#+��@{���r��ɟ��Dm��i���-"Uv���ۤ�Z����?�75*Ty�RЍ�q�X)0�-���b���ڨ�b�\��[a@�|�弄=�6�wA�g�6������/v]�a�M�S���҈����y=��~�1#�c����-g�|��R�(�Vw_0
�]�uv[���\N]�)������Fh�[W9�:�'�T��'�sČ�:W��<o�����ce�u[�S���~m�'��਋*�ԑ��1��o*˘�W���.o��! u�~8A7�� ��q�$�"T4	�H9av��(݆����᝴:�nSQ]�&��J>f��.�əe�y|�]y��rQE+/������Fk��x#�����ý1�/z�MV	�=[�f0Դ�ɫ'��Q |zd�p��`Fk	�Y��O�'�4!&X,;��ʬ���CĀg4�[A��:��6�c�N�6���s�m3,-�f��K]�#�<��3�7m�y�H}�����MH�2ӁK~�W��uO�C,2�[����G�S�vs�SD7��<�$V��LN�RG.�U2-s|3�/i'9|����"n Sٛ鮚-�Ǯ�9N�3ɖ�]0c��c���;0����r�Rx���W��� BYE�npQ��c9}u�<ўq}#�=��pO S�i�cϘ+�8&�+�h�e��P��]�\��ۦ�$�Ꭸ���2q�H���R���Q�A�́��g�G�xQ�g�F��UN	��&d�L�].���ۃQ-�qu��y9v� �
�C�@|��&�d& l@e��!���a�! ���7Y ���r�����h�p'0)���`�K�î��O��9����'x<�A�G����zu���2��˫����M����O��n���	��X������m�}�ڸX{O	{W��D���p;��Bgzsq�d ��ڍ�ץg1�Z���t�K%��qE=s�\N9�KhTZ�8�Ud������P�A�v�ڦo�&�AV����:��3}�_M.�sC��`22���y�\<&^j�q8��n,�z� �O<�e}޶�B�O�4g���g(4�T��5�PĨ��
l1���(��WK�o[^9��Ø��.��[�3M�ub9�����Gբ� -�DP��Q��b�2ʪD��Ն�A�N��:���4����K�'C�[)��(sY�WB7x����}q�Z��!�t���&v�����0�\mɸ�����]���*2)�#6���ԝ*v���T"8~#l���p��/�3��v��t�q����U.�9�X$Sb�\��,����r�g�ıoϝ�c3�$PO�tA�"khQ-�HAҼ9��u>m���J�9M�(%�i��e�e��[�C�����,ľ�(���y�)�\��d��_�B,V�Hs#k2�˂��������I��l��&/#+ןnd�l l0�^�m���R6�}@%4x�\�PLx�Jl�c���g5�|�Xҧ��}0�xrn=�>J�K1�֍�{	���I�=�#:]�7f�(�C�F�@{t$߸~�벫c�zMe,��L����*��R���&����l�}0�~��î�d��҄�������"��%�q�}bߔ��ocP��:���9�פث�*4Y��.&@�Fu�Gm��Ė%�-Y#F"�Eܺ�Ñ$��{����V����x�pR���
j�p���vB���D
�Ē����F@�ൡ�K���;'�y�J�.]Aa�}+���"��p[_i�G�'Q�с�=��,u*��������D��$v&�� f��%2F	-L���ԭ�8F
�l�̀�\h��p���i~]����ZB�����$5�ҷA&H�>��	���~L`n�ơ�q�1#�ChUqT��xa�q<#-�E6�r�$$�[��۶����{h||�|D��s�Z��@�G��b���y=�:%�9����u��T�%F��@�z�x����W�D8��u7b��S_�3��(϶iK]%�5ʋqU�tޚ�� 9m��[ȧM���C�Ɏ�� ��i�M��e/�
�����9��Ⱦ��pX�G0�m���>2�=[t@ �A��u�/|�D�]yPK+;�ks����nb/�3Dʒ�Eb�;��>p_���l[�-�f��e-�s����}�7���at�J��̥�A#� А 5��!4�4Ɨ�S�B1�a�6w�y4�|;)�Z�^2�F�8r��%�.�N�X"����ګ2����k |�}��.��gh��#���c>���+z��z �?�=���S�⥻�z0��R�9w��5�<lF���T�a��5�o\r� �&�>��UQyt�� �@2{UD�:�K���_��:oFXm��;J2%����n��:�`J��di&��[٪�����%���m*A�/Ҵr�/|�>�O���_�PJ椟z^��*���P�u�
!~������Gs]֜�Eq�ɤ��0w�Sg�j[�D��T��\�e4T�M������٦a])����_�s(��W�`9A��B��%�y�iNӕ݇�{p0��[�M�㊗Qڏ���NgJ2о
��̎�����t؜v��IrC�Hq\ǈ�=N�.���-n�K%�B��3���NC6��b���&zU<S���~����R��4_��c�7\N4����G�Ai}�6W�@�m1t i_��*�9�9�E��&�/���