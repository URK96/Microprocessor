XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:
���f�7`�(i5ﲻ"����$QP"�~c���~8�A��0�60-�O#�ɸ0m�JW�%q{a��7��D���̏�_=y�[��'`E�_g�U�Ք���Z5��E��|i� ]���!X>�h֐��������˷s�Y��g�6d+��JX<�` �af��vܐt!PЇrJS���|���P%�B
}-0ПP��E]%�\�\�5�w�e�8�����	���ʡ��� �z����h��݉�x4P)x �Ej���o0�����4�|��{2��N���QNY��;3�J�1R���DGA^v��#
����Mų�7��GT��� %2f�6����%*$i<�β�R�
�tW��>Z�ԑ�D�Y��@H@��P �翵j%��~�Y_ҨO������vr���Y+x�P\�9���eWC����ݝss��L���ǰ�ݨP�缧�gJ����k��d2f��0��Yf�'�}����i˄	OH�o\� ��K_��D�r}�V]?V{�	E��jp� $a�u�:���ىoJ�3!W�y�z՛�z�U���$8��ь��5��Y�I�1�:���S�̈��|�k#m��k����ZG7�!X�O^9r�t��K6�}�X�u����pm��3<�_U�����ph�>g ����̌f4�(��, ��-uӜ󮵬0�}�֯�|�����oG�f�FО�I�6�S��	f����/\��9-c�y���"C~[�i�/�mXlxVHYEB    5a4a     590��65��"ڡ���{c����#/*�M/����W�Ĉ*��/�>��kQ�H{V(�7�@��q��6�)�1ٓ_���.�>���ți�d��4C;;g��_�7�.Ƕ%%��:\��� A%i�h�X�Ɨ���wɬh�^�A������X�\�$��v�PL��x ����aW���Ch����/0x��0�IU��!�r��e/
���{W��@�����E_�V��zh�W�,T8ʷ���Fo��c`�eI�� ?a����a�����9Y��@��[:�iaU ��k��Y���z�s��:�ߛ���"��ʸ�ha�����ʲ�k����+��S�\ʶ�g�N&o��  �<����x��)Y�9�l��2"Ea����>á*��T�u=�u&�5��<��t���Ќ7�<V�F�Y^���u{��M��K�ɋ�5��������sn#��9곾ɭ-�B��V�,m|��:6T��}�؄�2Q�I�ܛhX���R���)d�Ye�pЖ�7g�������-�o|������=\�5�x7�h n�t9�]�Ť��q�)�)z>����k�~�}�D�#��_� .���M�r��[o��tfd�R� ��!E�׼�}6��!�X�r��3���Ӿ�WOB"� ��3�"���9�;�i��	N���Y�WnG���zs�,�O��vt��W������r��A�"�k7�[,4�5ڐ��E����B�K���p���?��D�)�|:��G@Q��@o{�C�15%<>�&���� ���Yo:T=-���}r&~�&�dD�7A���1���S~�f�����-ph:a�&��p��g{=��oI��������18_t5�,��@�_�
�$�ݻzcQ�ҏ�5���u�N��s9���.������qCl舰��%.=�<���3�Bg�c�'�4(�y��d�;��o���tO<����j���lT����j��zn"����x�z�n����q����1k9�����9�ڎ���=h�H�%t��"na?�@n׃L~�ܻ��GJ":f��6$���p�9T]EE�L]��C�r *�jU��
���,���3 �D�]�|I���B���CH�F��R@�ѐ��
��r������xg��ܕ���+D��]	��S��I�������Tf	��I�Bl},�G.=��<ќ���I�[D�Y �eU�4�(��+38�
Hg���Y�Y�É�T!������X��
{�:���W�C�����v"!�R��1hT�wr��ef&i������e��@:�����a�}�kª��]wT&��[PX[ws���&���h�";A�ߺ���\;�e��z^��S�-��]]n�j����  �