XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3�b����]Amoc��>_3�TE�5~
]|�v6x:W�O�c`G>j��aC�<Ϩ�K� l���!z�d�����ve:��/�۲���O���f8��e�U����B�@�!��������a.�����}
�rm@#�����'�q�>��}Z���WY���WɓU�Č���?�i�/O��#W�	zE��I��s��ɹm~���`BI�J��-��sA»�]X��h{s(���p������*l��#δ����;K/ʄR�V���A��p��,���^��;TSGҰ�|���!!`��P��)��lOk;�]'���޻"W�x���r�+���)#���	+�'������'d��h��L��b*�ɳ��
4�'�/����F/�z�:�����H�׭��=�+�P����T��ٶ�@�|�?����(��~��_��z�Ӟ:����TZ��H�1��Zp�l�m��eC
��S�Td]Я�S /Ǹ��X҄�+n�I��cE�����i	6l��Ak������G�B�j[�����b{��64mI5� �C��̯��	@��GfM:y�Ҵ&�b�-��u�%�,T���V?=m��'-�l�E%WK\NS��쵁�WQN%`�*)�K��%��u��+��]v*��ŰC��_���2_���4f�w�b�����Hw|���'���?�d�G����mA�P9�		d��O1����"`����!e�۽БGklgM��,;b�F�� L��s%�XlxVHYEB    5ff4    1040���K�j���{�����L�LNF�'���|M�
��42�˫AM��h��nzt�VP�e
u3�s��Qy�v���R�l.�^i�	��7���$S�vh	����j����r�,f_��	?�>P�p�gs8���_l�9z+��m��������'.����RP��6�LqA�Q"����ع�����Ti��h�����]�Z�*�I�Ch�\l�)�&湇��Ҙw�����[�=��Ʀx�i㬙k�uߵ�割e\�$��Dw��W���b�܇��s��J��'.����>HLx!D¬�,�_s
�12c�`�  >_��Fm8�|�VŜj�\z
��!3^�8BR~�hU�K	]R&��c�<�2���%!�y��-��=��{���m 'QB׫䷹\����T��7Cu�0V����\��irR��P0���-�ÛN �l��:3��iB��qU�/\�˨��/�58ey/�w	��$�M�}M����Dϭ�:��e���:h����ǲ�;|7ŵ��z����Z�P��FJ�mٽ��Zr�k^솈��^o�I��D�#X��o�\�U]�O�zY���<a��/w<l�'�tm�0*�_ �&+ Y3�!g�[l1^+�T��'�'NOB�KU�|�땑���-7�_�둪�̩�u�9$�Q��%�s27�[���l��Vy���T��O`~K "��E��+~���k��ʯ�D�_�~L�����/b*(Meݖ���6�����cm�7W�0h���9���if��ʉg:���и	磧�U��A��ȡ�m�~����h��}Y�n`�.E�hm����"���-z���s�qcB�s�#�&8����&p5�$���CD�r��蟗ZĨC� ���Ĭ傲�	����=���Nn@S�bG��e�d�L36��a�x������j��윃yPZ%���>-'�N(�FQu1F�)��!�@��3g�0��Nͮ34VO��r%_s
A���] x٥g��Miw�^�JEkmkF��est��ݵj6�Y�|�/QY�1�4؃7�ѓ�6j��������)FDX��Z&xQ+{0B�2�qCN��n�*EzX��[��Q�Y�>äB/��NOO���O�MzG�� <��'B5�O��~�u��}��G&"pL�r� JΫ틇��Z�V
W�FUv���Ңo���7)�WYg�~v�j�J�#=bNrf��":P�`��(eUe�\�P�&D��܄��~��u>����*�
:\��v����mR��nWC������MK��&T�4RV<��OmZ��?q�X��;�iZ�,���4�.�h����z޵Xﮣ)�T��C�G��S[s��IЙ�*[��f�6�I3Ϩ�9�oRI��WT� 5eIg�Y�"����k|_U ���<KZ�?o��ᆑ���OU����9?�0BI���p+C��r�����1� ����)H�͹}�78)��{.1*���W���w����Ew��}����}3K�+��;�,�.l@ޫ�:kC΀�ߖݕG��A6��q��ޓ�l�:?��j�
�$���ƣ4��D���o8��k�w��W�������3���SR�//�x�A�O!���IXҧ�^�q��+<�c�w�JKl$���ĝ~愸&gA��&� ���2[P�!��1�65T�[(�X� F�ξ���Թ�8���,tyi����Ϟ k=o��7e*V�v#RSzH,�T��@�F��=�m�m�c!����'ٔk�wS�_�^�i�}�s�@ؗY�Zu�r�e�b&Rg2�i_�s�dϱ�_%Oo�t(��Ї�pL�-� �r���K3��eAaT���5�4�Ѻ+O�l#Dwg'�S��Ə�s�b&�q�h/w��Q�m��FN���i2��*]������}�1�!�;�l��%�k��m%e���	73]HvQ	B�.�+����n[�`:X�x�3��mqR�YW��nSa��p�V�ͷ���� ���d���[F��@���ld�['�%�(!r�yh��x�ʧK��^���_��B(4�5_!�����:�i���Ͷ��¨ft���Ъ
��^7����21ڑM�P�R�̋o7�|��%Muh[��+�m����x]����[������eS��z�Dt��4�wf�%�lV��y��ϸq��6�W�&u���_h�:�_J�- V�	̿�B@��w�i���݋�F��u;4��pZz�r��{K����9a��Q��s���uũg�<K-� �.��ɜ�G�)O)��bk��E�bZΣ�������"��E�eo]���M����N��z:�Q�U��DL�t�{�]�8�1��X�K���J^m�+é���3�U~�4k�u�=ڿ$�k��n|�*���@;!�'{���a�
1�n������A(�n�ڷ;��hQ-�մ&h1��`��i���'3/��T�����ov�*�B��i���o/�A��LW;Ve��{��~�q9Ӊ&�bJ��2��8orз�˽��T�z^�l-�m	!<����Y]���({ z�ثׁ�A�iC,��~���<�h�b�n.��#��+��`�qF�	���;rDƷ�@�2BW����\����`�+����!��ꌤn�&���g=D�Y��Q���3v|�U���2�H�E߽�,^����Ϗv�O�b��Q{�D��D�6�1_�?���3���`��'�EƼ�v:'�ԙZ:��'����S�9x��w��K�c|��t��HȮ'�˺�!s��q�ʹל���x�篌�Թ.���X���p�� ����̴!�Y때�E2�#�ZʂL�E� bn���va���]�p��U�ڄ4:��(j���Q�z̝�-�ƒ<�`?}�����_�����ж��4o�Y�<�JDT_F���D�?��j�r�S`7��R
��c!0�n�I����^:���8O�#ڧ��$�oЊZ'cA�#��Y{�*�&�5����}O��0���~[�ŉR��mpX��4�$2p�����S�N�W����,on���i��6[��9�gH�ڡw~��9?6���>ZWL=V���4g�֍�v�t�aoc��|�+� ����Ft�]�����HMlJT�AG����E-��N��(-�i��{��̦/S�F�=q|�[	�9K1�$����d�N����I�.�K��^�O�U�J��QD�'@y�Cm��U���WbΥ<�h�E"<��b��f6��\�?�He��ֳ]%z���I��q^
è `\z��~2���W�=/RG��+F�@Oh�U�����cG6��
|��� |��D�۹g�C,D����%*�{���;����qH�p��-/��+��ٌq��wKP#�d6C�����	o=!�&��I -٘S�O3l[����쾻�8�|�X�
*�� �y��))����E�=�;{\/� ���K3���2�P����2�gʉ��֣-~�[uy#2i����g9�=�L���=��W��_�[*��?��pLm���"N��� X
C�"��,?���a�nb �*�l�N�Q�-�f���g�n�0�Ы��y��b�7�,u�����{�au8��� _����K)��Uђ<� ��(Y�ĖY�"U���z�3�o ��)�9 Ӄc�a1���W\�w�B�C�@$|/O�� ˳F��]��/
pCܠ�z5���M�)�i$z�6w~�"j�>�;kVz�����'�0�R�@*H[����)���j�]��☼��wX`�qYO��1����:���e�9۪�e
s��@Gr-�/�e���Z4d����&���.*8�rM�ڤ_�e���j�ܳ:Q^!��_�MI#���i�K-k%f ��c'}�]@_���&�/:M��'j'�����{�p#�i�������
�N+88м*��c��0+�D>H���Ĺ��%$ܢ��ʡ���Rp{�P"mygbĻnC��ql#�A��)Ɖ�nW��_�& �
Be�a�"�c@������+�1��WPJBƙ���(}]��_nݍ�K<��سh�UX 2��� Ε��+_�F�