XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���M0
���T��U�f���-{�;����M��9u��k���e��R9,]	k�Dl�a�������?�="�<�m��;A�[r�UD_*m�� ��FG�o��;�}��l�# _��{}T�283�z�f�����s6�d�	�.]�2��r"`�n��KtI��[
�K���M��g�[7�v��Mћ<�
~O�Q5�ϒ�ԡɱ��a��O��EC̗I�
2�Sn��Zx�� ��g������/���	�����Ƹrω�vnpC��Ź�IH�rȰ�Vj�j�0VIڝx��+Hv3K:���Պj�/N�3�d���@��ME�EW��
�n�\����v�}���4�*�hQů��Hڼ��*cy��^NS���ќ��,xj��,�%gX�6��\��%J��O��0�#m�åZ�f�?H|L?��}6t/Xެ��)c&��(*ꄮ�I��a�M§-VI T ��9�XC�ΏiOAЯ���i�eÀ]��h�@q��w�ę�7�{�0OU�8K��9M!�w8�KW�a�Y^����~�pe85��R�����a���4{���Z^�����I;
4^7sGgG��,�n�W�G	���y�=��D�&�_Y0o�'+��o�2�4��J�X�Ԝ �4AƔ#m2L��AXH�(�œW�3�Ԝ�*��� l�ї��������O��T�ԩƨ��;�ZQ�G��6E�Ka�ak/&-�Q�eI7Z��c��o��%1^�-<���HXlxVHYEB     b35     3d0­{c�������&�x'{�i�*
^�7�F��B����ʖ}�$�QSE���yjo���z13�s
l]�(_@��y5p	�ʢ�΋��v� �ה�L%^I���_O��4��+9^6�#v_z��?���?��Vg�tӹv��gR���	c"`x��ǭ���~E�M�Ŏ"��E�Sx0�o�3O�C���]��|x���w�-���V�'�͠��ie�Bxj�?�q��0����Z��1�H^�A�5�tQ^6
	T���� N=�����J�kM����:�R-�z��<o�݁*Gr��oq�Ȉð�I���q:S�з��Z���0�>ڿ�g�Tjr�=p�%�5�un�$/�w�g����w1V��hQW��A�����a��:gDʂ��q><��+��I��5t��Η!���w�l����YO��;���+y�ාt�B�J�ŲP(�'��^�⏪�6�DU��-՛�AV6)s����4�`/'�=������Re_��U,2����}�)���A9����Ν%�������TlꎉdR6���4���O�@��R��)��}�xA�p�'W�]QISx�����8��rx��3�^1�jq��Wv�� a.(G"��T�Jh?Qn���
�.% ���YX�^�k�}�%��n��N��F.c��Uav�ISD[?�KI� c���b�� P�E��s3��f��!�Lk5����W��k�5��՚+))��d{��+���#^ �$�BDvC�={|���VT��8����Q2~�Mק���9���8�a�g�YTI�s�(S΃��r_�0
I�A 佾L�`urXq8�i�q�e���5���2��ئ-�s�!$�+�=Y�z�;�r��(:5�����b��?�8�xOs%��T�L�������q�A�^�F��s��2��Y�WD�7�Ɂ �Yg9����v�"��{���X��ن
��