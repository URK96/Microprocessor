XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����%���+�R1(�v0��͖:s��R+�Fb�]���8���6�o-^�̯�tT����f����U��pt��>�X�9��$�q�K�{��ʜ�BRn
���=ֽ��,�p�l/*��C=r�I���>F�Oq~���Ͳ�*N;����(P&�O�A|��4��.[��$�0F����� {��Qɤ�.̌pNc��Z�5�DH檒�>(s�A��@g?�$4���'H�y��VGP��	4��@���c�1������X�@�U�"܂�8�r���T%nf���#���T�^7�[���;�w�_}y��- xz;k&��:�Vv��&M���FJ��\��I\�T b�DAA8��X��M�b|<�4�#�;˥�t0w��
��S�R�A0]6]*�S.���fK�`�qA'��M�ſ�M$��\�aB��89�7w κ���M$S�o�Ynk��n��8�t��0Jv��.]l��+��-�a[�����O6)l�Y
re�t���z�}�`�K��찔�@�ެ��<�-�%�۱V��U��҉=T G�k�m���϶�1e�30�3���2�+)��#�ҁM��:Bp��*�U���݄�����ʣ�t�ڷ8�O� �)�ظ�5�����T�����Q_/�j1h:fX����V<6j��Y+��Hi�� Wj}��]t�Š���4R2�f�^DbS�LM��ڶ�Z��e�q���g�l���zQl��{��Qs�?��=�!6���"XlxVHYEB    7a0a     c10���~lw����R��E��mC�n�J���{ݜ�q7�Q�^P�m+$�����x�I��2L3�"/K}�_)�T��e�ˍ溞 Ȍ	2��7_��#s�%$h���U>���=� �u�>p��=J'��&}}�v�m�8zS��Nl���ͺp����uC�/m�i�2vVU4wd�JS3a��ک�z�4�����:Ѐ�<em��2�-�>互+l�ٲ������<b`��B��xP�Ƌ��nm/�"��(F��)Z=�NŬ��GP�k��!�c(����CQQ��(7�U���K�V�=�)�`��g����"��x;��%�,[������IZ3, ���P��xq)�h�/�������ꎃ6�;U�a�A��v4(�L��,x`^��wf����f!���Z�w�t� v�q�}�HT�v�Nb@�2�*�������	�x ��/f�f�k��y�N�%��0�wߡ�T	�ܓz�j�ž� ��E���>�,%�����d���Pm`��U[�N"�.�E��:Þ	����؄�y4������1˨ե��n�h�bWq\�|^p���^�ѷp�/��,��i������˒��M����V-t�<&Re_�3Z?fށNF����?�(,S�š�sp ���U�l� ����0ubEg����J���
�$1�Ŕͯ�t?���	����[�S���G$�'_D{�pø�
��=��;����kv,:T�>�X��u:�����s{�T��E���	ٸ��|�ȥ��F!l�Mu:w�֤�u��i_Σ��CLH|�b	>���n�n;���ƣ�TUE��}�T�w�x�H]p�̡���J�#��|�N�$5��F��:ĥ�3�s�?GpD�&�O�׭�zX�S�e�Q��������3k��p��rS�4��?�n/7��9�[6�	+r��tV�(��C�Oπ.	� ����H<QO������*�Ė�t��A"Q^L�e$T�ҿ���^YɆ��`ٓo�F��c �X����L%��+���S���a�Ѥű�恚m>�v�"��/H_f�����&+������GC��P��DR	W�U�@j�sP)�m�c;D�NPC
�s!��V<kU���!���6�}HkA��lk����q��fNI�{�u�f�������Db��xr������|Zw!�����NU*-`$/�ӗ�.��Í�T7�a5u�O�s���i���<\s�t���.��&Z���fe@�(���Mp̵	��KB��v#�<`.�o�T��͆C�괋�~Sj�~v5鑈4�j�&Ŝ��� ���2OH={K��b�3�>��\:��K\��y;��¨h��׆�Y�&PG:�]�ZB��"�Nŧ��s����͙��*D��D��7~�z�I�gԆ�O���$�<�W�O ����Į��9	1a�O���|��h�R�<���.i��Q`<�����:c.թ�H�䏺�E� k��p��+z����F�-3X�Ĥ���m?��v�_��]���8t7(��hw��0v��>]��P�0 E<�.�E��`��5�������[��+����ٻ�<�,aޅ�Q��*Q&Kd���c����������W��L��_wHti�?���)
$�h�qk�����F�y@�9J�gN���X��V�e��4�zm���EmS�Ag��!�u��iU1�8�3p��y��c������&� ����?���Г+#�- ��&Qm�x�&�hMKg�#��3į��f8w�"�g�Y؏�O�e�<�@|���$p��ϔHoɰ^�t[e��ϦY��{�r���
�?*�In5&4��dv�YLю�iE �~��Jbڍy�ˢ̘mEwn+9�r׫M���>�K��h��$Zڣ@���D<������sO]}���FȆ��׏.��v1��2�
C��lK��Rm��<�";~`�n'Y~u�I��ǩ-�f���� Fd]ۙ����8_R�X���F��=���`�(;T@O�NX�ve(�nphIO�:��m@$v
�Ň{ݾ��gG^Տ�O�/ �dF��:u9���E\�,g�nq
د�Ŭ*�}8(D"�#���������a�^�Z�N\#&I+�g�S���²�����m	���HK���hko����M�j�k�2.`
���p<�wŸ4��_�b�R���`W:kSH�}�K��������5b�$�Q����fv�#�"�G)�g�i�W[���X� �[�)�rn�6L��_�_�+8$\J��11����8b65+��X��21�ġ��ʣc�+	�쓭�\��Ө��犮�ɫ� �E�bE��[̫k&!��x7c�u��΅I���DbH`Y�VK,�Xq��Ư��
;�L��&�%@��Xܽ1�H�[���Ih���iBAt���T`�1,B-Q����L��᱋���t}˝È\�8�:E!���e��x�;*�P��Y\ҙb�o�I��e�$��F�%W+��R�#�ZRZ���	ي���{I[dk�|A� N�y�j�Ě ������d噌%v������~t����F3�j��ԫ�m
h�VyJP8�����Nv�!���V �]�����U����Xmݔ�h����Ά�9�+�VJO]`��x�m�pv��+�Ja�x�+Dۋ;r��B���؋����祩&9S�D�K��}�C��Р5m�/:�?����ꃝ#G��osl�μ�O@��0ѕ�)$�	m�b�d}ir8Ke�`�3 w�+-����[� �9Z��yN&��`����t ��~��
�I���;km�U��O]�&���g�������)�:~`�DU�p\An��v���Z�V�GFT�#D�	�u����� �4�"Irȸ�}�G�:�-iT<C�6�INg��Ձ��$���E�u�$��׏֡�S�+�z�#$J�A�a��4�5��2�}6�Sz��ݑ0�l�E��.�3]!+~nc!��
(���q��j� n����i"���3CuW�1�S��`p ��=w9��C�