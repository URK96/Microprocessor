XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~��]�)�R&֫����.��;0AڭC��_��{�7�Z�g��y�:{�E��x�&��\�����=?ѭh8C]@Q7cr�w����Z�1~V@K������֮֡@AM�"88B�d�Fwu�w��Үqk��p���3�,��7*�U�m�g�!�����ǁ���Ktv	Owskjldl�b_
�k��p����+�q]��<���Q�!����� ƋI�Dܲ@�"�.���X�3�e�%F��;a�z=s��s�E���۬"пW�i�Kÿp������f�QB�^D"	U�F�W���N��<)���\����0��|��W�3��Y�tm�3"/6�a���6��7U��h��\�� ��g���]��16Ƈ�`���l��!��Ӹ|�7�&����LfR��2}L����1Q�>�����P��`�a��W霺 {tR#����7KR;�b����<D�Nh��b��7w]&�6%�:��Ҡ�s�V@�x�e���Pr�5�!x����;�J9�Zq@CE�U��������M��~C���W�3��� �C_�A�m��&�W�v�tcz���g�%��Mn"�*�W<�5��ET�C��H���-RAѶ��lj�%1zh"��,H�k��K��]���0�.����u���iW��)X:�A�`�o]��w�M4��h����aӣ�گ��#���c7���j�v�׶�l���?��䒹��:
��>J� 5�z�cMIa�31H��F"Ir��\���EXlxVHYEB     935     3e0�o3��v��L�o�;}���*v���� ��4�;�i�p���a�q���6�{��>�aQ\��yt�;)ʺ;*!��g���B��v������h�!�$������~�Cچ�������NK��Gw��X�|_iܬ��׆��Q�^���������=G^�l'F ���J�YŶt�o�U�ڵ^f폺�6m��g��+0W�O�@�YV���ɸ�z}=*����vN	EY��cQȇ��@��V���'h��A�ٺp���=��~�eR뤂�@'��n9�S}kA%^��P	٦������𢯦����.�zϚ8۷W4O�x�w�p}W��96?�|`��QתJ�!��PhX��?QSMJ��sqd�\̣�����(��u�^�����
� &wE^7T+7��Ç[[ic���nX`c?j���NzئDgϔ�ʄ{��:{kW2���LFE�)R�g���"���"�n�ы���_�ȫ���4V	=W���Z�hN_�Z�nF�]�*ѷ�Wa�6�k���1.?�ZЬ��6�/G��&���o����-���{]�;�>�@<��4����b=������A"26�� ʃ0�;w�K���^v�N���K
����)��
��Wώ$��]_rz�R:fE
>��������گ�^�AN�wq�<�8�e���(�.O���'�D=�:���0���H�ߥ��m�9@��2A��'�M�G>S�;�b)���	ר�,t0 <���N�/�;�}gA��Wg������N}���p���dJso�&����E[S�s��ֲ���������!�hN
wN�)g�v~�\���I8�%+���CO��K9�_��B�K���LI0�Y���Jн:7'��lOk� $.�{	��2&�"��Y��r+���R��*y���$Fv%e��GQ���K���!r��]��Y�U��=�F��t_C��Ĺ�P�t�������$