XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���I@���4{�l�0��|�����rh���?o�:Z�$�vQ�6���t�Řhޚ�W�]��`���wT��h�!��{ 1�b����b����:g���xs�g���~oxǵ�_��E�N�w����EI�]���ZK�ދO�.l��cS���x�>��@�Z҃y��R`9B�.��;��j��p�
D�ApFm�Ͳ'���P^-��u�܁����@Gl`M�2���vB\�V�����i&,{4��
��c������QB��˶c��s�����6��>��[o��O�&�*ot~п����׮@+�u=[.�H����������2���'A2)?�IWo~Щ��a����4��H5�co]I�	\Qp��r��Ys����M���Y-6���6}YM7\�(��ߤM1Q#��y�N`�Ѱ�<l��d�{a+&{1?�K&pM�����p�
�Px�g��V`0�<�a�L0h��x͡��'m]���q��(��OF�1~h�d��!�,��{�n�Cr�a�2"�T���0X6��Ae7��/��h[�m���6J�$Gδ������-�Y��nct�h!AH~��r��⿇�yH���3�	���R��Q0�$¼Q,.j�t��!@	W����Ϟ:�W uL����W�]�.�L%At�q�	+od��n�eɁl�3����il@��qy�[�O�l�>q_��e)�H�{IX�H*�x�꘠�pUWS"��]����	`�7j�<lXlxVHYEB    7e17     de0 >'Nt�򀿋��$�o����z@�So����6���#���%𹅷
*���'#�RY��_��EB3���)Q�� �
}���(����ș.]d}�s)�'}�������U=�I�IuYџ��M	7z���M� ��څA)�E�BRR&Z�u��Q�f�p�%�Y�\�Y��mc?x}�Lb韭N�r���vu�ګ��tVR��<�K��� ]p-I�@~`�a�����l��S��H�Uo��4��kI���\����G�c"�\�U��l�?��-�B!E$�/$�r59�Mj� חuh?��/����3y�ւE|?!�~���#��64�
�g�C��������Lwxvȴ�-K�������JŢ�'\���ZpV%�n��I�#!rǐxE�Rid,3�Ш�3�*��q{!�yb�n_��ӭ��q�f� 'Q��+C��p�u����|�	l�l�&��H������s5�eJ�7ԈnC��V���cＵq�\��Y��F���2W��=))�ny?_���u��A��������f����$�j��k�l��h��T�U#[�ޚ��r��AK>�1~pɔ2�[����J�r�S�u���S��p��EC,�~�+��{���dM%�*ev�bT�����@/OC��u��&7/O̜LʔтI4�Y#�b�O���Ԥx�!o�hW���(�]}/v.)�b}3"�Ӈ�!�EX�yXo���\r&�,(��wgl �=GQ�����nʵk�����(�4~y��IjX�$k�O�0�w� =G����E���}���6O�J�P�BڦH���|d� ֤H2�*���AF�Ő{��F�qq�F: �|a��,`�^N��6��Z��!0B�ϵ���)��`��k�!��u�	?�ý���x��:�F0rF���#"��a�*x�Z�N(�,z	Ȇ$�i��+��~��KO5%�����-G3B������]w�`�,(��_�������-y�
���`�U����6Sv2�ґңy�L��"Dۭ�}Esݪ����p{D��s��i-�:�iZ��3?�Jz
�6�DU���lݲ % �9{�Δ��rJ�_�
��R1��z+���t˟Ɵ��yXw�Ԁ1���1�
���L;�v#���G|��R[��4�o%F~/h6FM�}�vߨ,��n^����	�P�mz���FI�K�~���Z��`�ܙ'�Q�8:*Յx#e�u��C���W�xwء�U{w9�K��)�c�V�;�9�,����Gs�xA��]�N{�lQCc��T��i��u�&�rINc�R��[1��ĸ�nJ�m������H�˥���:F��z%�ǩڬ7�h�j���.�h�%����׍HP����%�4�BTy����8�y�}���u�Vh���) w ��k2��B������V������5/�dqr�&��]�a,b�#��X+T���X�<���"��C���&N[���S���+_�$�E�P������i���nu�w��.��yغ"�'��b�q�A�aޤ�x!��d�t6i8^+��s��>{�r��j_�|��PZ0}�z$��α`��nXb�ߴ8G���~{rKNĲ��Bs��Br>Tos����W�Ee!7mI�5G������-�[bW�ɾ�
]|ͬ�ɻ�W��B��S^U��=�Out����6DhQ�/�3[�4g��wAk�.����U�nA������zV@�\�"�|'�����੣�%נ��FA-�&�u�_�>(���BT�4eG���#��S��oE6��h�yB���H�k�s��4�c�A�0����nuz޼K�����?�8la��1l�~>h7[x�)�՘� 6�����Y䑿ó4�GZ0n1��^�����'Q�I��%J�s3�Vv�Ŭ>����䞓O�}?p�	��c����L�O�r옊W�)Xc�f����Z�4|/֫d�@�� �n	���s���|~���=R5b�:�7F�5+�<���ʮ�4����K�ׅ��zM*2�-Rw�����_E.x��^�D�pW�����$7.� !!��%6�1gS���	��S��w!��UB&�i7
���4�-�Ɨ^�V�1���T������]��ڒ�n}K�Bܠ+�l��Y[!��'��v��A�9��tV��� y$��n�[��� ���U\{��H���9)��;ȗo��%�3�!t��	�EL�����,^2 iDy�р���|��I���쭾=X+�oR��[�M��2����zRe-��Qy��V1���x�`l��c:k�QL�2�0j����S8�<T����Z�5�({&M����0�6���I}�&x�z�ɒJ��u6��{���S��b6�׫�һP��ԧ�F��7�k�y�� ��~�1��O��*�SM�{鯨�rq��L��5t���Y�}7�Th���p�VY����p׋3��sc@67i\��J�3�O$��A>�Hsi����lA��u�;�z�GЛ��n�;��gd��Çol��+ L�p��<�ײ�1�R5�a��V6���?���b�X�%�jKW�W3�@��&���&�iq=aMř��G荷�_^��E�#�ߝ*bC�*�*�pS"\T��I�L��>���$���v��3&��Z�zcx���\�7��=��	��6�<^{��cS�9'�7�����K��hŠ�TT���]4� 'g��G�
)D��+ǟ�y��^ G~�S��W9��e��i���D;�_[0ũ��PHo��9Ÿ���;� jpQC���@`�W�?K�G
�>pY��n(�}wH����4��=����a�h��P�'�+|��c�E�i@��ѵ��rm�_<q@�n�p�Հ�����X��; ��H5G(�'�GQ��<<��T����?�+,E��UvjCw$��>,;���Zku����uVZ�d^(�ӳ^mSC���F%����u��$e�
��X{s!���l�=|͍�g*��$\�+�����ˇ�@���8� /�m3�D�U��Y�|��5g���<X�69�3�LQ�G�sO���q°�i��H}��$ZD��Nܻ�Q��ƾ��,��`��@��n���q�<J��ȐDw��b�w���Ws�vvVnI-XY�v�@R���ꌈF�u���L)I-��"\,�tz��R��O#蒯���J����T�A�a��س��]�Qs��;�^�\�9�:-�֬�/���6p{�${�q�:���V�
��L��Y5� �H��\�%bO���O,���[�"������.����*���'z��|�r2~2��=������,䆫]+�0��\U��c���������8�,�2GG�X(@���%��>��2�~8q��J��2�l{�⊶ES>/�&�!�xf�@o����l��0�T�^	�D����#r��I��n�vLr��R �<EY�����k�ql�E|8yڠ����1.oG�,�BM,Y����SS�yT