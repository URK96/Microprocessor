XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���߰���T ��Q��ǡ��0�-��0V*	�{@�͇�FC����*�|����Bty��H�ok����ȯ�~����Ь��Ձ��Y��~�4ߴ�����eD��.ٙZ�	�C��<���� &����3d���K�_�ne��pX 溅,�������󢖄E.�w
x����|#�q�w���W���s����]w��F��'��Gl�⡓��Ӹk�i\�=/�e���G����뭇���W��0b�(%I�1�g��J��6���Keѱ�`���3b���M��j3�U��N(7�2�'�{�@	G���wZ�a_f/����4�(eZ+��܌��R�Z����B ���ߪ�s�B��M���sL����!9&h�.�¾�!,p�L��$�q�8�h�8��@<r��Z�2(�h���n�nV��f��y*�>���H�N���y,Ԯӱ����Y�Dz��ꁛ��l�n�ْ�[d��v�3�1���q@dA�/�S����D����W�*j>��,	#���J��ң4�����ɖ͊MNF�pѳ�7c��T�"�'
��^�����Gjy `}%_ff��KY߳w��ӟ����Q+�Ji�%�3��WV�s��sQ�z�'N_��]�ѿ%�Hc٭!a��Y����o �=,�&3?�a�k*oNh̗��\k�_�O���L��\��U�-&�&J��G��Ix�|�i��'+��m����5:]��ѵ�����������a�XlxVHYEB     82a     300���[�?�Υ�x�UŠD���'�?"���������r��q倆��L��?�*���[�Y3e���Y�p�U�1��\/�&T52t�$Ao���3�����(,�w�m�k�V����v�T�ۘQ= �|1��>}i$�Ƀ�XkJ#�nՈ���SK�5V	s>1!�L��
�}_k��G@D��VĢ���A�Ħ��?��*)�49��ηB��DP�X3j�K�fR�T�>삉3���?x���`�ͧt�o�L��;~3ߌ���
�D
x��n����rv�ߗ 潙�)���q���ӚS�������ვJ����N��㏭Q��M�oߵ?������nxȬ�EY���M�j�����
5�� ���/��C�ޞ�����k��'M��3�l��$I�)�v�u�N�"�.Ɩ!k\)U!�	�P�E��1mw{��B�}���M-O��p�K5�Ϫ�=_���ˋm8�����*݇�Sc(��ʤ��	3�o7�����ԕ�^�.3�Rse��\en1�c��f��	f*	��Z����e�d*/\�jk�����"�%;�('B���B��l��6�8X�Jdy�����j�����C�2k�L����
�c<��H��	��̆\ ��CIvL�]��3��-��J����}�S�b�K{w�=��o����)�U5Wa=^)�{�|L�xBO��Q�z��[��UC���Ӆ��g��	�Ý�?��ܳ�����Y���}����ϖ3��~R