XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9��D�`k�K3W�K�gT-�jCE���v�H/��~�"�B!��Dfk�)�h�N�Hn�!Bqθ�^���>���u��簃e��\k-V�����Li��w&"�4�ڟԗ���{n��?�������_)Kjx���^YX���,���L���h#|	�5$9�&.��&-6.�5�mk"F�6�RQ\V�g��}��w̢zR���0G*�����(���h��ЪMi����[=����Q�GI"�� `����*��.�K�~��4���+"07,���.ͩ�N���I�ց�7����/���+�Gq��+>�x����Pߠqv�s�� �z7�������Z �#��̔@.�ض���16����h6|0q��XE��U���E�D���vϫ�0L�䶘&�����Gd!��i����2���y£ԏz�7@K�E�ɿ@PX�ؖ#�1�,j�$�I!��hPm0�MV	��NE��� |kK��s�d��(}�2��r��i3k��N�+�М2.��5��svB]�w�:n�%[����5��j�9�3�4O��!qǒīؕ�!�A)��gH��P"<�5�]��l@afF�bK>g%�ZHj�ϟi����?3MA�1-��]�Z#HT"~�p�c>,�/#���z�	�cGy Kp�����Y���%�b �Z�J��x-5�V�~�M����	�
L�~ihQ��#(�߃W �"�D	����y��r�|aI�R�n>�\��5kn!�XlxVHYEB    5ff4    1040֣u�z������k��g��yYIQ�i�+~��=�`�=#K�2E�b>֣NTk�;����u��X{a�E�s�Q�y��Y�7�'9A��x�`h*0p�~P���1�'��-#�t�wS������T��{���Q��yWע[�K�� i�?�y�Av8�����3���~Vng�X#?PyGZ]�ah�]�����8rϧhh�pX��C[�Z�*�Mjn�<M��q�׿�	�+���~����L���3<�j{t������-�xl�k*[	�n9�\�C'Ɛ��eV3�F���~�C�X�O�HY���*�&#���;5����Ք���?���A������p�ü�Z�z,?f�����m����E��ou���qj�ې#��*�$I&��9��x�����n��)�����O��D���l ��-�X��_~����V��P>���N%�	-*w�%�l�����9��נ�X;5$ �E��p�\�
E�yl�p\gҁ	L���hx	h�qz��Y � �ռ���|s���h�J�;�>��S��$�-�YG9+�Q_���ې'����<�0qs��1�}�$m1�5Y4����]�,��RȐ�|I��IH����r)Q���������7$��OWc����6�h�6@̩�7rtn������y[��*���� ���#���3� iF!�)��(h0�v�"ʹ�
�3SB��p�A��8�D@u�Z�%�:E�=AgYX�4�Kj���|fp�)4�HΗ��5C s���um-�ݽAe����St���3BE@� �K�I��
j�
�;�����}�bz��3�_>��o�6����7��IN�?L)X]s�N`Qj��G��\�-1�����H@��<V�{ؒ�a��]�dr���^^Z�%M�I	����$��릍�+�b���b�]0�Q�T]fp0	ԇƇ�Bf��A��T00��
{TBܐ��k�X>T���nQ�]$�?�2�=SLkS�˲��eE��7e�Ͽ������zM�ao$�r�ʓ�WA�=qyyb�J�X�'g~�Nrp���{q�3d������M7-橠�&R���y2�D�f�C�'6�����7��쯭W�F����i4K���.���>}�8�ۻ� ��D��J�ë�3�2\���?�>`%����Z~K���6I��h O&�>b��lS��Xjr��
ю��������0#^L�xEJm���_%��L!������ԓ�*�2����+���p}�+<�mQ��<�l:,��޼E;�#k�g��T�˺�}5L�v�C; �@)`�mG�/�z@��r�t����4��H�MA���aq�6ܜ��������l	h��1�u�86���a��i߅/��EEߞ:� !�K�w�n�G�T�'��2cM0��<-��=�w���s	wj�a�E�` �䁒0�,�7n�
ݾ�-����Fq��^�CP�BR��^��P�D���+LY��A.y��V�]l3cڗ��[͊s9bk#���,+S�K�����vu���.¤���N������l_72?��/�9�%����]8+K�N�BcSX�qCf��ɞ�0���3�o�M;&���>��ڷ�	����1�/]��Ɂѯ���lz~z����Jn���4̩�P��3��~7����N�f�V�����o(3"ע�ze:e`p�[�E���e`X.�Y.D31��h֟=�Q:�J,�^���5�Z:l gI�k&���d���T*�&AhM�r�}Ra�l������"-,�FgP[F�iB�,�n����.{Ȇ�h��.�����]#�c�73gj����[�<���54�m4��{>t����P�yB�1"�3����V4I�ΆaEy������ٱ�&:��لZe���ȯ?���Z1��)�%����z"��n�~(���y݇@�>��S��򱴝�A=|#����}��C�ҁ]-��[�M���e �_�B�[:#g��?�C�� ���UZN�-���S�	��g�K�c$�rmL,PƏ?��2:�
T���gϮ{��81�YzJ":��Wh���q@�=+��bY$1F\�4�4�v`G#�hr��ǝ�vFY�0��pX��6�}a��O?_��)-�T���M��U��'Dx~���;��˾�٭NZA��p�����Ƕ��w��<f�R�W#���a@`	�й���H�q���ķ?-�kh�R�`�u�.�q�����n���z���#�s�>��K�T��g4e�:lYs�9�U'�ޑ�^�G��9.~v~��>�l���-v�
/	rI�-{�Xg^� 
���ӡ�����g��C�W�]H�p`k��1�I?=%�{���i����;r^�t���E��9t�А�E{�/DDh����4Yy_l{mtB��O�
��$d@�HG1ix��p2��-��ˀP���oEN֙���-F��醱����~�Ǌ�t�}U����{o
�"�d;�Ķ��՛EN?�ܗ̏`A��iǅ-��nbC���>'��Qo�l��:���m��P~9�Һ��a׹9;NNa-`��S��:�&#jE��ee���J��\�m��ծ�,�+�8�So�>��p�d�'�jq@��f��pS�#f�d�_@��'�� �Ɛ=PnM�q�}ͧ��m� r4�!I�6��'�"�;��l�Ǟ���u�S��E빙��3Z����i_�B{�R�?�N��񉔢���|#աq�61:J9	AÈ�O��A���O;�pn7~R�[�~LR�qw�ߑicEX�Yrk�¼T��v����PX�Ľ{r��-�%��@��s�����=0�;��[Fma��<i$C�j�*��F�_���jY0d�C�缇9~���W�ul��d��ܽՒ8�K+���������k���y�^���
�4�#���So��j���da��	s5Q����H��KS��c��kKB���8a1ω���� �I�+�@���9C�u?tI{i��^X͈�~ =p�>=��t#�$LcQej$�A1-���RA�9L��%q|e,�'�-��=�G����!(�sՄ�B�+4;��*��j�ra����w����5(���D�0��g�רּ�A�n݀��u>��:g%9����j��5�d���@y�s�R��8hu�W7�C�歊���r�p����9,.��Ka��������0�1X��󨿢{	QN'�O�����
���m��#�oS/�(�y�c-$�� R]�咊1+=�x�2:�����R��(f��BV���Pf�_�r�|AL���?��F��Va-��t�F����E�4�)�\�\�ɕ�I0�V��]M��_D��/��\`�Z@�`�>��Y�>S�x⑂�<���O`�MS��ʒ�6Z���ʋby�SHd�&M�oÀ�t�8a/��	��a�jm3�ӧ�r��/�����PÅl/��>
՜Y2i~ܘ8M��E&�:��t�7��Q��ݻ�U�z�Cb��f��T^UԶHfRUv�PD�V�H$L`�fQr�a��:��7��RP���A���G��a�i�vx�T�٣����`�~���A���œR{F��tg��	���[?Q���W�x�#�y��
*P����	��`�&�(� �# /0#�����x9�����8!�{'��n��%������RǱ��C<-|����XJD���nEp�A�t��Փ�(�
_�
����?���jc+�g��n�.W|��V��Q��c�y���ߌ������ f1 6n3.c�A(AG��EQ (��q6u퟊�)��K�#���_N������O	h��0��!;\�Ȳӳb�����!sGLn�����3(w�C�@��^Ț#�g�����S�?�8�D+.�s�5h£����g���/L˚�"�|��J���}�(qL6���F�Uw-�Vp�z��x?����f7�`w��͊*ƨXi��n�!�G��������#��;�������Eaԅ���a�r͇k�\0����H;+��Z�U��6�*���yS��q��	��$�,0�~��~�	