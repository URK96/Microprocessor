XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&��L�E���-��l9F�F�@hD(������vb����s�AM-�ܟ��z��t���>Q�``�6�te��rQ�l�8��(�J20v�~�:��pԧ6Qǣ4r8ʱh� 7b5����U�Ϝ��*��6��j��:%�2*��]ᡷfgtM=1?{�z�\J�}�8v<�k�~�����|v�I�qBQr��V��rm`:u�"~�д�m�RN�녚E��8I��b���=�0��ts�
�Њ(p���7���J�'�TÓu�k�?8@�e�Ah�����^6�p�cK�DQ��axv�&��_��rQO=�>�闩��.�1�s��|�pohbW.D�%k��bQy�ܩ�$�q3�x}��H=�_���~G�0]7o�x��&_�)�qqF���J(��8q*u ݠ�H�2�].��M��ض�R���N_�-����i[O���xE�{�ص�G�Bb:���8���`�/8-�jV�pø=2��<�~�~~te��x�D��ٮ�8�V�>E���~����̝i B�8�@UXg�E;$2e ���c�N�>�H��A5B�7(��i��P�T�W��W�/��h߸h�jc������t޳�&�c�M��ε�Z�H�:�k�_X�v��)�Z}�����-�[��=���X�г�%�I9̞XH��Ye���(�25�"�Q�"�g���׭Ц̾և���,�Ģ�j8�m�qX�`��{�ܡ4�O�9.Ƴ:qq������;����9�����XlxVHYEB    152e     580���sԨ�2��KZ��o��v��jF�#��KX�v&%�oV�/�9v�?A�"�u]/{6�T7��ن B�b��9�����5g��20�?�;����IW�um��6? ��8�;�+��g�ԅ�￳����� yˡ�O<C�U����j��;��#E�D9��uq�ϭ,�\���ɝ� O�p�xE4�75u4���Jn�s7U�W!����lK���8��X����jg��
!ӟS���}��'$�R�(r���pj��)u+�w)��"��0�36�)%�+{�ưG�|�ʱ{�pzR�I����ŋ1��J'�;�mX���9cg2IL��]��(?�{�q���	�����w�,��8O�t������h��	c� 7��7dB����y�q�"v;�kή.;�n�)^m������*!��4f��^*�h���7+��X`����F��Y�,P���\	�����^(q�aP��q���G�3�փ�Fb��mJH%�m�>�7b�sU�|9�U�Re���;ճ)�#Tj��^E����Mݡ�<��.l�?�Kݲ�?,�C�Ǘ��w(����z"Ė]�e+ +b�?���ߟu��ψ��T�5��t����ka�OV0�;�9MM�ؼ�aq������Z_�#P��o���m�͆����:�
^F�;m%�m1&�s�΁��z1�k���t����|_�wu��5D���?Y(6�,;�F�CK8�G��H�d�j�����(���HC��y�S@&�cӫ�ϩpltI��W��_�	R�P/f�v(��{����5�fs%3�Z��{�i��se�ύ���Y�j�y֖KM�F���HYu�P:�%��Lat��>t���_m �*a�w�=BI?����p;'�5�C�ꭒ�!=(�R�cG{���{�������bX!5fN*�*ltE	�E��[��=F�ڭ�C]f�If�kg:��Q�xcԂ֌�Ģ"dq�����?��V@�7uM�JZ�s�bW�m�\p��c�� �T�ro'_J�sZ���9*�`�S�C||H����bϟf_�\0_���d����ZB��Z޸ٞY�m�bj������G�?��/D�I�.�D��LJf6������E[3�������_��1˴j6�d8�������Ϩ��Rt�5|L�悸A1n˓�I۬g��nK����	 ���^��߼M���L����=��B�J��p�݅@/`@�yݳ�W�`ֆ����-!/���L�%����?�@:�[+3D��+�[>8�
�����G�\�Y����>Ey>�G�1c���pD��a��� U">�����)��X#(_'���BS�4�<����/�u/�"���GНFaoq���ȯk'n	8F