XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ڀ��] )�l�����VL~�׉��ھ��@q	-�Kj�񹦱�y�NWTY�bx��R$7��~Yg���X�i�b�x/��m�y��㓘D0�i\c�:��.i��W���7;�c?qbؘh9p�Mv���-9h���gV���p�+-�m���+4��D핯�L�ba*�69����?'�� ��E
�;b���s"7Ёxlճ�~�& �S	K¶��S�)��2������8��h;�`�a	ۦ�h�i�~QFE@��-��`R8	�uE���1���s��݊�+��)=�(�B<)�X�^���a���?/�vv�[�	��s�%�5-���[N>r�j�7�Զ�hH���!�Z�[�߲��6��]���
W6
�ď�'0�ۤ�ܜs���w�t��o{.����������U��d�?-��0�-!O��_*O�%��g����9��OGFV���NAPD�]^�>f������}�=��o�9H~0K7���!���u�eR��3��w����������?Gi���w����`���b>CQ�U� ���m��٨�9n�h��g�6�w##z���Ȱ�Vڤ2w�b���r��Ҿt*�"�Gx��G��9�^/�,�6��%��7y��X�㮁z����k"u|�~�Kf���+ITS�}��P# ���f�O=*���QX��b�jR�|�ԛ����w��R��CJf�o��GՖ���Z��A�h���'E�t�"kGD��O����?XlxVHYEB    1cf5     790okEͨm�y\4��������Λ"�K�_9_�1�y����>�UB!�S�hY/��Y������o��L
���:��(طkgD"�E�����ߝ��Z��<P��}kH�k{�t�&ԇD��� GYF� 8�J6Ж�X��P:F����(Z.,�D�����F&]�g��{ �pX���WK��Ս�b��t�a�͕�`�d���A�_��=~���=���}Du�&jVy���4��VI���5B0ㆩ|�G� ���e�b@�W�t�d�;A��^F���.���������$��L�3:��|�'-�/+i,��x��E]��z2�on~�K�{�����u�ȑq�A��V?�6rv`Dӏ�rP���ȏ����
�?�5�k��{bY�Ӓs-�# E���jQ�ӯ�S�n`��������6=0ii	a�&Z�ex�RvGE��ik���;<��=�x��ڪE�C��:����ƌ\솢�$���֫�c�Ru���A��*�g#2�M��Զ�̈n:<�i/��)W�����ךM�` tPFc��2EV��Ȇh�u��ȁ��}�*^0=�
�u\�)a�r�=9I�YXP��/'�k��KLw�a����O���҉G_�c��ν�yM �(5����F�4OӢ�۟�����˗"�B����+wt��'&�
�.Z��K�. ]�Z�2���"�No��z��T�I����db�.K�p��e��	�&������#���*j�cT;P��y��j����:<�иc�8�fw��0dA�m��9��#���Q��$�lUZ�<��ٸi�z��=���,n{�b ,�8��&�B`�ξ;A����gS����qpH,
-g/����N���q��I�9}�Q�R�v���P��=����^���K���-�eE����h�J	ѻ2e&d��|-H�A�P�#��v�A=�Fso�����-;�4�vQ�W��{��.flS�}M��#xI���J?Ǹz���3�i�՝����)<!s? u�m��V+�@dK����)C'9!�+b�U&�I�ٴ.R��?��
g�z��k2�j/�ň��w]ٍ��f�7C�i|�(n��%��P�`COY�L"ڧl���T��1�xc�����X����E���jZ: ��m�O����B�T� ���Vx��Z��"	^o"����_�	Z
��G���@cW�q>�R���$
7&��k�x(�q�[�[�UX1s�{�2%fn�VP`w���Nx/���e��
���Ɂs�� %�p��\�h�A�,K��D�ѐȉI�����2��ʥs5�[�5NMڹ�Z�J��Az���/p���LS�V7� �ϲ�~�ZƑ��a?�����e����� ��#7	��{3���'�A:E��i���c8�Oh���&�V�)z�%��BT�C+o�&8��jR�T��&�p������?���﹉n\-�e�Vx��%FG�5,><�� a�L�50� �$�RxP�n/﷔��6ϯЗl������f��P����n��R;`��\2�\��&�G�+�\֛�����|����f����\� �uS�ֆ2� ����s�^O�\��~��Dg�f�5�E�𗱂FB����*
����;!t~�!N��*cM*��	lp�0bs���%
7sDhi��W=hZ,76(c1�;=�%l�L�v�t>&�����/�3]�0Mq�x�Tg��{j]���bAf�Il�t�ނ�$�&��%��e��N���?�+��ַ���xŢ?�C
�+�;W	v�F؎�Gha����z�H�����*��e����n��d��J�$�nk��`�.�L���;I�������\�*�di�	�S�߉*B_(ڄX��oi ؆S�9���ýqzn�薵P9U�N@��t��Q�y��J�4&