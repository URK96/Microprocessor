XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����zK�á��6�ZYx�������T�4�2�F��B'���B�`�
��E�p\�ﱧ���Rjeߍ7a	������>kP��:��SߐDX4*��"��f쉎���{.�;���x��tl'�խz~�|���=�huRe�����g9)Dc�V��x���Wt
P��5�)E����C�*�ԣ��A;I̕�4�}n2�e�:��?���GCلy�����C�^3]"�kzW�-5��"��m���_��_կDC����_��ֹ�G���gW��f��U�C8^.�p+=f �k��_���_JB���P_]���:\#�:��.����0�>^�46� 0Bc�qp~��i=~E4S�T�z"kpV>�"FrV�!bA��P�')+y�5���� `�7�*e�����cQ��'Wʰ@6����
b#�Nt�A�VL�u֓�o���+�GgP��8)2�i�:�p�?8v��k�J�g9&8h5��t�<���(%�<�0!����k��_vi�b���E�q�c:l�˃��B�7~�7����Ů���J<y(���v'`A��0�`�[�P �����'?y�/`@i�v���a+��q]��$�%݁�R3Ͼݣ$
�%Ѓ5��P�U�Ԡr��벢��2�N�d^��\��F�Z�������U�m(���ڸ���K�$'7���1�w�'�¢}�~W���N���,*<�gA ��?)l�!�g5̱D>�o5OBj�#�����b�{���EӔc���E�AZ�XlxVHYEB    26ec     8e0c�d����Y����1-���R�-�4υc��Ư5�ڦ����e�,���3&��bl��O;�fa�n���d�-9��&���]�V�$�a"���C�=�H�J��#̱����u3�������sgJ�����GP�V��ӂT�s���*�֑��E�fZ�`L��>�;ʥ�5u����X����gl��F�~���n���_��˃�K��Cs��a�����@ǀ2-�#��)�~�ӛ�o�����)^�����I����&���ٱ;E��e�x*3�^���j	n����.�_�À�G�yp5|��}�͐�N��y����i�aUw�s_�v�Qk�/o}n! ������nݴ|��QN����� ŏ���}������.H>���@S씠�U���J��īW��6��-�։�����'_����o�zH�v�=g��;Pu2�a�=鸵7i37r�
���=�[��^Nܸ���4��?ҒH�Q�T\��?����JX7��|���D�� P���{5�S�~:�0�d����KIB��+1�C���K�N�u� M\��R��m\�힦��N�)�vn�"�wL�gr��Zt�uIs��2ja�j��Y���K,�LV�&�o�6�w�C�~`Mvv���߰4�&J��r+�P,�B�.!h�>�H*����#�zC�'7U�Vc�5�Gs�*�4S��e�H�9�W�O��,,��{u��Q��:��acCt�,|f�M�%�
�p}�AY�m)5��?�.g��)�O��gZ7,'�V�(�,$�I0j�\� ��\��M
�4s��6i;���_a������4�&'��5AmV��AZx�\�W��!��jɧI�����2�m��ZI���;p�}~D�b��qY	�}>LQā"3���(oT"k��L�@"�+�k�wנ�YD}Y����#r���l�i���/b���1C)u=���*�	�V��g�B�a�O���t��O��T�C�O����h���1Dz��qRbb��V�^�2�Y�m�Y�<+�� |8�q۩�T�f��2����zL���$�a�����,�1[����;���O���3BC"��Z���u���:f��8������;�)7�'��<���������O�2ts� O}�	-��]!o'�dxV��A��V�W����s��V�C2�2Lab5�	�I�n��j�62w�ܲ`#�$�P�w�ʿ�URtsu��xw�%r��:Ɍ��̈́b�(	�� D��`�x;~�:�z��	�*���%ä��Fh۠ɏ�mZ.��~�e����_F	*v�u3��>(-h/?(F
�E��Bz�5Q�J��!@e��aq�thC��I6�׳�V%j-`�qOb������A�H��6G>3�m���������n#�'^��Xy�����o�G��8�ˍ����8 {��U��k拉y:�A�Ӌ�mF��'���"�9�͊� *^M@w(?�g�Z�M��m���2��� N��a?�Mڹ���m8������">�?�nܒ��V���ƿa�?BĦ���q"��<.�䚬�So�w����ӇF����Z_�]]D�	���������.�Ψ���V��X�o�	H�~��
"ayC?!�U6�{>�%�դdl�����wZ�ʭ������+���KA�0`"�d2��2�6��s��a6b���@�}u�yV��n|�cR�<�p4a�j��=� �=�OQ��^Q��S����A�B�� �Ԝ;9�g�~A��&�#��.�C�e�Y��cr
�2t0�Yi�'�1��f����-M�<p"���ձF���͍������_չ\�h���$B�]MR�Jۯ�F�c/6��,�=����w��U����#��̴-{�&FX,J�6c����lZW�����QLM��`|��6��Vg�|d���o�*_���Q�wBGn�` ��^�oT:��n8����/4�����Fp��g�4RJ��%ŔAR.�>4�)�����wG;HqsC���E�k ��Y]ʏ��M�>Zֱ�r$H�?	Z��6g2j��"��M{޾�r���f������jtǑ6K�s7�M��)�� ��V(HN��ِq��{�c_ ��
�Đ}(�~L{�٢������z������dv�I)7;���D��vޤp��I���J�k-��a8#ɦ\���U8w����T�F����dv��H�W��~F�