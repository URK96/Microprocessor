XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���d����ǝM�ֱ������w%��WYa��k���T�	m�G��o!o\��xY Ϭ���0���D�8=�JW�]i��:NpMZ�����ʴ�C���G�����DD����5�<k�H�N�]о�jǌ����+ �>�*@o�({�'=)��RC ��T�$�'g}\N��Pv�@�X�@(髐z�&������t��~ei {,��H����r�^+p��E��p�4�5�'���B>.ƕJ�-"x�+N�\��n"���&�a�������V3����	�߼��3K��[%�~��lb�Dѷ�SL��~�d ��uZ E�1�)�5��⇮�ϱ@��Y�K�9��e��ѹ$~ހ���Q$d�+��+����N�p�tf������ք�J�7�>/�s�x�Q#�H�8F>��ʨ,\�c���;\��4�u�0�߇l��؛��@���3��2%]��V�[,W�aR�K�f'�cޏ�Ed6��qd�r�t���� �U�
2���E�ε#1��Z�V��� 677�r<���>��m����y���{d6/�Q�뒙��I��"����6u���z5��D��p��9�vST��GktoGjJ�UPP� ��S̱�����;�Z�5��[���nR1�ڒ�#[�@�*��J�B%������q:� �'��8��3x�!0�prp��)�8�(0.ؔC���_�Z��ae�Ǿ!C^����	�Qw�7���"�;�RYEMi��]���E0(@��0�XlxVHYEB    27ed     8d0C���ge4y���Q�o|Jt6�M�wl=,�9.�˰A�J�1�{�j߳bG��5`���<'��p����6��M�k5b�m��yT`n��fT�C��Ǟ�;��6ѱ�"�#��o�w�(�?���;���#�?Tn�b�n��My]���Jv��j=�;�˼���9Cf�&�.�fCA&C�Q��b!MLX��9��S�冽h�~=d����#�����&ymg<!��m˗�h�V��e�t�����ŉ��2��3�Ѭ��Q�ґ흨8)�G?��g�K��PȻ)C�Ԟ�3�H������#x�g�����̣�*�=ˇD`�g`!K<5'%����&�=PK8V���W츢�/L��fЮ���!�}Gi��î� g�L8L���?��(N��z��1(�8ү���z2��\F{�Hd3j��Isf�fWn|���b������T)b��s2�q�7H���.�����v��ֿw�7�H�t����9�^V$�g�hC�n�ךS�&F�8&��PT)k�����y�M�6�I Y"��	�0!�iR!,Y�_������d����\]w�ʩ�
��4��O�޼рD��t~~��Ք���������
a\�q�Ny��� ��};�=���.���LL����Oy��	�P�ϝ�^������
���x�⥩鉘�Ls{�O6|��fk�>���\<,�G��c
t���0^s@ZC���PJ�ll�L�_[,��>g�L���Y�����N�J�o�ƒ �ي�0Ϊ'�qł�� `�]�,m�c���.L��,������$*��4�0�j+�/"�w�*���VULe�P�H����v�J�æ��|!%�GB7y��;�X>�D)W�9Y�1��s����u|;���-�K�M�����Gf4�=���H-��?��N�`޺��l���G�y��R��W��=�6_�v�0/:���̛zy� =�vZ��L� ��/\c�&Ak���HsJ�B_>�(EV������3�����x�-P��,K[`M3�u�{���o{,�ﯓ֨�N�q�0v�E�i
����O�G�xfB$���S�V��j�7��^}3�)2�5����ے�d.���5�@�+H�����6��x�v��)����|���)��� \�ڟ��ĝ��O땹�����,8������E�O����ZP�&rQkC�x��1�>�:����������[�qR�4������{��*E_���ƾ�8�`&�p��'ۂ�4+���Z}A��r@6ce�oc^�p��z����C���4<�Ā.L��8:j	��'�l?�HO�aämA���K��/�U�IȬ�ϯ=� ��_m۠ˍn5��6����H�d˯���[��l���%b�n���p�'MZ�(ܭVC���:bW~d\������~\�믭�.e��X++h��ƍb[nX�P�bɧ�t>�0�2I�'�gTܭ��U7��U i�.l�&f��`�.�!|������+�M�v�h�����"�ظX�q��i�G�7�e�Ŗ�=�  F��P�{�{�;���_�w�C�uIY�󰮞��ȁ����f�& "*��J	��9hx�G@��0 B�9�G��-D������>��:Hg#R
q̎Bt�G��Oz�y�αΠ��"��M|�s�1��^Q�����<�n߇}Zy<��ƽ�Z���;�v�� bB;N�/���Jc����w����S��Q`�ˤq�Y��r�Y��=�B  ��d�E�^�6�D`@C}{����������X�^r숌�M2�N�����L���1���#%�LZ��I�5��?�OW�.��K��yi&���5��uy�D��u:BI
E�����A�6t��V#yj낫��_Fm��m�����hAԁ��*B��㚲M��,�T5L��|���jC�,_��^�t�_T�Q�%eƇ�o�(n�iG(�u�!���OR-T��'[�|1�v-,�~bB�J�o�%���9v-���^��9A΄\�5���DQ�q�z��i�q �b�S��}��wU�8 @�&.s�b�C/L�0�=`�]ܚ@瀇bD�E0H�˭����6\�� �}����K&�O}��һk�u
q����sx�~D3������AsR;��<�#���ο����΅P?"�+UZW�.!�Ω-K���j}1U�j� (��X��ҕ)����k�;