XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��őe�3�E���t�-ř���%�I���@Mm(O9��e�-�Gg��5���W�C� L	R�e�Z*��%kUJ;���狞��U�[r���5aQ�:�����N���q�p諑���䩑-.�A��b��^G�����H�h	���J��7�8|�W�D5M�P�˦��;��1��?��x��o�X���NSw��_"i�&j,K��kM0�Xz}<3��a�jk���z��k�l� BN��Չ��] ?谤���l{�i���a�6�Vxn�a�d-.H�S��2���^Y���Y
9��`��?s;.��tc�!��X7o2�'����/=Ne�E0>&�p ����8�����=H�U&b�t�t$B���L�+uP��Á�!���}*�� ��#������(W�;���;��!w�l�y��P��>���tr���8d$YB��{3GS�&A=�g��a2��h&��H:˹s�K�3E��@������� ����qmNSOX��Q�Ϭ�p��9��yq�=愤�,J|Y�{�'�	5�Y�~�˷� X'0�pJ�i�)˿��"t���y���>���3ǢZ�ժ��5��F�� ��u��?;�Q�\��mokN�ۗ�R"d"��2t�E�m��W�9&��P��0o6;���J+���(��)���-ًOtz����d,�m�v�]Q�q�Yi��z_4����o&_�_��,¾��:���-��6���`P�f�a�5s 97�Jix&�B�~$��Δ�"�#XlxVHYEB    15c3     780���qh�Ӿ|j����S�K���i�Մ�!�Z��6�Fxܮ�p(h�Ձ��^x�`��� �>���\�x�&~��)��'�s����g^�G��&�u)��خ'll�Lf�:.�@A*@�g4�[y���,�C���W����*���cE�MX]�|ʞ�c#�E�{�M�+�˸��Z�QӺ����/�#��N8�VW�c0ǥ�̲e�V�&�E)>:-#=��ܥ��0�-��c�w�:oe��;,E*�߯��.ݐz�8�����H�FE�����	�n�ˊ�Wx�7`���Z���^�4��Ms^#+p�b���g�g+�.���֕~7���ʾ;�|<O��Z�&-��.�|bH��|O�)@�B>Ҏ�0�?=���4�Ic�<�篅���g��)y)Y�U 8����2	�0��u��)��#�[��4�,N�k1�5L�����u��WQ<7Y�>?��ih�_u2���)O����j�t������}� :]"*.��lǿ~XR�\��	��)��[�D����)!w�ps��:B��������tv���]��J���z����Ť0؊�+��Q�f�`-y�����+%Xq����P[ [���\��['?��o�~�ti��V�H+wN������	0���3��MB�DG/Sξ,7���IbǬ�R뗼��uG�o�^o���U�P��ط�V?��`	x=�� �M� 	���C��r�� �|�4�����5�Vf���m�#Ȩ��V�M�[��y���Z2@����D̷��:\T�W�q�蝈�!�1��E�a�,-�Q�g2\�VK+"��ҩ�E,��\
~�/���F��
��A*"f6:}
h��8"�yBߥ�>cZ��R�ga[�� �C�Sռі�w:��������1a��FRJ�78�:7���-o��%?����oo�������'Aw��;5�'�]��&�zm�xo�����L�n!��.����@�T���������"h���yU�R�T��!e���4d�U�DK,i(�^ Z??<s��1��7
R���,!�x�3��~�Wa�^��}��8�~�:"����h��a������7�Z���A�!��i}�n�r ����uD��-���K�mb�z6���ph&�L��1U�&�;Y=�r�5��+��K$��9
�[�@����TU���(�Ѱ�N��}>�Ī��#`�}r4��@��c��X䔕F����sOB�*M@�6�1Hv@�M��^5i�%t ���'q�깹�ŏ�w�?R'P���ٗ`�;.mx��1�`0��S�/.��h�G�37�7s������E� ���uT�J�7���p��Vx_�pV[Er(���տg���A~)	�Q�W"$������� ���y�[�}��.�q����np<^��RT.f�S�)`6r�L��߅np�F؄\(�0{�|��	<�w��=���]��%l�q�ĄF&����>��h���}��N�mobo7��ɶ؊�2c�WOl	I�F�w��Z2(D�'P�5n����lY���@�Y�Xg�����
h�G40h<͹�k�@�:4MA�����wʊ$����y�\�1��`v��=����E�>���ۯh�T_};���iSUK��T�(>��k ֨7�ӯ8��h��	�ƅ_� ��{��r}DV�R�_��ǽ[82(~��rV�0ǥDi�<�^A� W7A�%��"�)����A��,���S����(��)�ˮ�I��G���}z���	>ƞB≟�)�����%�-j�gi�9�@|�� ��r!صO���C9�E<�CVff����}��N���m��}�Vj�|x�O����y4��W�m�=C0�L