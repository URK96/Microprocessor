XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����"�,��d������t�����b�U)�f��s��<�~ ���OOk=� ��,?�P�eI�o�W�b}�j��/*�l��%;� xEo]�ͫ���j��P"�`�������Bj������>�*%��_�E�дZ8�p���*=��
�]V��\�C��na���(�t�T��9l�]h�R�^�b����\{��u>���mm���[.����i����wA3�0T2`�XJ�^����'!�2\�؏N��k���>ݞX���!��q��Cq\�2��dS���uL��M�|S���'i���JVv)��#�><��xs��Y�	؞�u	5�d�$��D�5��̓%ܦ�G<��y��MpҪ���X)3�sr�(8�.֗�@p	$)�+8�<���t�����d]��f���YvD���i�cix�I����;p'V�AN���]�H�ː�?㠜��,�#�8�ҮJ���ũ��{=�d��Ď���������p�{5��6��(t=�ǯSR,vD!Ф��x�@h���+��28Y�
�u0 _*�^i$(�ʝ�K�G=â��4�w�xt��Ȓ@��l�m-���l�}��B\[��a���X��.`�	�o�>-r��R�5,Qz����k��1�>�a�O���;���5:ι��V>)�g��%��yi�ѿ��D�E�}o�
I����H�X�^�Ԟ���>:1=��k��������vgY�?߱`!k�9��h}�0?�Ot�XlxVHYEB     b08     3c0/>I�=O�Ƣ�0�\i�edq�v�z����e%����cfß�Ǳ���R	6+��U����0��?Ƴ�\�P@8�xOgm��Eq>Z=����A[��%4Q���Sŭ�c1�]�rY[ZtR'l���O�^p����}U�I�a��wدV�q�X��@ZP�_@� ������ߺ������;=AP�e����)���d�eâ/g{T��q9L��1jV�>ԩ�)i�
"�;�+eJ�_�7r8��d\������=�c�H�&HWf$�3��vֶ����T�K��J?�<�8.]��JgÞ	5�&W�����EHѽ����p&q\�3"��w�C���Q�?-&]�&D���U���ݪ��ƣ�*����+����Z$��GY;��{�j�h��������멺�dFyp��9wKxȓ%S+�1.� H�T/�w��{8�>^�����^�W���WT��^���n�g�9��c��}�#{�J�Ȭd��Xw�It�8QL���tU����9���?�^aӮؗ�vh��j2K���J "���C�a���b���⅃�2��Y��o
��
��8���<p�fw
{� ]Ϳ�/�y�L�u؅�Ã��� /*;T�,�ω2�S�%������6��"��wr�D,6�V������K���w"9��p��c(CUfᒒ�V�Yn�I	-�x�mع2"0������S��D����5RA����{ᴛ�����A��\r��6G.˿N-���^�4��n2>(���#G��d�7D,ش��苆52b��eO��PKD�u(_�є�S��ժ>B(/��r>��1%S%�u)��Ev�e��Ȝ�@���Z��A����yN}ϥ5���Z��	rΑ���G�8>�j7�B�uܡ�����¥��ڮ��X��Bq?�� �FZ�w�5���=�*=^��G;��鉙��#|vyf�;