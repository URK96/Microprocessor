XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t�̘P����葻J¿��w��rVPp�*���kE��$�%:�
_�S��K>W�J�(�:�ܱ��SN~R.����q����=w{F��i:S�v��0��9���Vl�d\��h�²6iRW�P� ���y~����ϗ(L-X���`�E���7�\�n꾯����ڵ�k�P^�PG
�{�k��T�T�	��P�M@���P�[B7x��{��.��J�3�ے�W>��0[�<$�9	����i��7�*6u�*b�R.}��aZ�Xu>x�w�ؔgߺ���q0��4&��+��h�3@�KO���8&�D��[�x�n\j%�EE[�w���|���4_?�h|��ͅZ
�9���LE�co#���C��Or�(+DZ�p���� &M@ck��%��-P����RЩu�h�.�;\�f5R,��׸W�{�߫��.^ �m+���+��"zY]`ۻs�G1U�h�Ψޡʄ�M*f�"-���AҬo�����U�Dsh/�;	.ٱ��z�v}��e�.Ӭ�Z@N=Ü�%�EV�6�`e.����e7�?�"�uH8~<�¶I������Sf�z/�N���n%2V\PY�����}�A�*<6?���zOoC;�<�g�����J��{;�0*)Epl��t��G�Ө�2S��S9�Z0`�+~P�9�#S�됶:X�N=-av>�cX2Y�������"0�����W�c���#	X�(���q��}f�iP/��8��.��dz�2XlxVHYEB    1585     5b0���	�w*�����)�%��˫URs6R[�m�8mux7!Rqgb�I�M������q/1Q_�<�T����Y�������ƛ�r0��A��-��q*R�TԸ/'�z��OM��f�b�%�����Fr��jtĊ}��ͻb/0t�KL�O�ng�Y��J�k�¿�?�F��n���6��R	�q�����"Nۛ�˪U3�D�a��XKo�5�ñ����L�1��tJ<B"�Q��%<����n���1j���9�O�
��vCe7�j�O�#ޑU�*���:).�3띎H�ن{�n5�*�� �������Z�������e�9o��0���T��G�(-봋�&��Ճǽ���(�����*2��|�'~i�� �?00C���N����8���l�H&��hhN��I=�K�^��Q�����xs�U��zs��"
��(����z��E���F|"�ݠR�����#��Q{5tگ�^(���T]88�A�V7L�-P�*���ˆeh/r;D�R������?��LU����+��J��jp� <��X��=X�k]]��;��Kn$ۙ�J�������n/�p��L��Vҭ�9B����4I8��o=�&�wSmLY�YN׫�0���*���?�]I��pǘ���T�$ǖއ	�{��Vذ���s�_��ű!�.$�,W�7�3�4�H�2uP����?�K,5
s�*���8,�ګ�������̓q������,f�Xc�L�A!��7�H��z�Mg׶P�:�#���9�w��j����2��;�cR��Oi���I��=�6�~T-�rJ���!/ιC?�]�-+�*M6��-�����:X��FP}ΨFa���zdu˘wa��x5�-5#��l�t�RzBŻ���Z�G���z�9�g�VxB��}(�i[���"y;;��O��y��0�kGI�MRlZ��~�a��a�Q�}�����O��C~]Y�J���IӍ��=�k����M����F�gcw F4��A��p�+g�4;�V)/L3�u�!�S��r؄s�b�a +�Z�e_�8q�;~�'������"�(��k�� D��|0�j#��M�U�����C���Y�,�v{?�(��S��͜��-̷SJ�9��[�@L�����$�N��=��u!��<��G����-l��T��j��pHP� |�h��)S�QV�%��a�8kRG_�Nj����T,ZNe�nD�T��g{k�7�dB��[	�OwNW�������/��� ��<k���ĤH�'^�Ch�b�5���jH�	C�tq,����^~Ny�j޸v�o��t#��ָ���\��6��~>�����E}��T��U%���q��T6"W�a���~thΫPcS�c��֦xX.2_��!<�.B�U[��2��
�嫧 M7�\�<5