XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ڦ�J	���@�$��3�H��!@�՟��rN�h�0�p���j��+�3��+9�+�^D��|�L���s>ޛF)�z���e��١B��&҄b���ϋ�z��7�$~~�jr����>&��t�)m�Zt�Rh0�Ii�.3�ʎ٠�Z��K/�N+�Y���O��$����w��'�(�v���*Yj�g8O�JJ{��/M�Ҿ�8�[�����!� p�0�˖����7b[�k�c�p�N~m�=@k��&y���/4з6k�]���t_�Ĺ��	�0`7�xr{��F�5Y8</�L;�Q?��|��$���q���6~o��� �4ˋ=C�
��3��bh�7�c<�q�;ʑ�V��zd���֗���m�pw&2)X�65g��:Cࢮ� ��Ͷe��ȲZ��,N�c���K� ym���A}�H;\v���v�/|J����S�bZ���zW"����y��No�<:���w�\�D�3��5��=�@QwR���7xq������t���j���'���d`�+��@.�ui�L5��G�P��3t//��z����ڱ�L�a,D����)�q���^�Ew'w�$��PI�������;u��2�9���g�t��Ѩ=�6����-i��M����S��zW����7V�uea�ĭ�]�U�;����(6ҫgˋ:V��.�:e��)�	L�kʉC��\�n;R<Wʔ���ZO��u���H��G���m2� @�N�~����XlxVHYEB    7738     790���d��p� G}�
D���e�,7�$�n�/@W��ҭ�#�Er�x�{x'�aƄ�)�x��8�c�~`)�=6Y�;�B �{�:C�,�p.6���;�)�W��z��k���σf�Ny�/��R��^W�B#��{QB?Z��n6\��@ua����w��>��jbV
�<�%��|T ��?�t��@�(�VlZQ�x���;v�44�K���%�8(�U7���X�Y�r�h�U�̢�r{E4��޴5 X��f����󷅽�!��S�cs|�Hɤ-�����DX���U�ϭ{�߉�K:�z�B�n_Gf�D�U���v���] ���5�u�!L�`��<���f	}��U�P�$�ڛû:�TѼu���{�3Ҧ�ظjQ
��'6$�Uk������"	�n�0�}�{�ÏQ�?kSjInR�3��C�~~-/s� ZnaͿuw)P�ƣ��@�+ax��A4l5�rz���T���P���aV[���s+�[��\۾�{���|y#.Ĝ�R���U���ՠs���t�"�۾򻡈uo@��+e1���}lJi}Rbx;�O�ц]u@�9o!֞�^�^�9�j 5>1ڹ�c:�%l�s�d���X��'�ɕ�8����2�����3ɺ�(�t������L���QN���[cë�Y��y7���Xe��\P�U�=��ʋ���.o��a�����<R/��^���P�U1K)���g��f��r����<]I��rB����1�����������oz��a�����Jٷ��N�}M6MV	����}.��S�'aY�4�M+�9����Y�/ �d!����Ս�s`���=*���~�bX�շrJ>�_'���I�ç��}W:�])&i�o�����=��|���fWF\����:Yz{C-� 
�~���8|�1��-�O+_թ���0�|Y���N����p&վ�L��hY{s������|�z�f�9T�ID�&8~Ŏ3 e��|�JBT0�^�:�p�_�$�xr�W�Cy�w���M���qi�FGxd	ܦC��\j0�U�F)�^e��D.�)4�����`��C�.�g���I{ju��7�=�����ˤ� S�FVJ�+F�զb���9P����ܑE���M�ʞQ��^@��8�"L���<�#�~lQn��#{�G������"�OyV�rV:�[��/�lH�H>KӅY�a֮�-l=��b�6����w��K7(|��\R�!���c��+�U��m&鴯�T�W%�%�׻��v�~�b��9�Bx1SDY�Gh�b�)�,c0T|��u@�q?ۚQ�༘�����W���lޡ�XӮEv@�.���]!�l�Y������s�I�KY/�\�����eM[�krV����[��Im��M�rU@w0���鿈��1&{Vd1Z�-NN��ې�<���58үۭ�_��C����nok���܊`�̸壽`?b\U��IՄ-f�:�j�h��v�����"���V�?�Ǡ�s�V_Wvz��M��Y"�����Y<�	��<v�f�!��a�v/iއn�D��(Wۓ�&���o�B|p���Ȃ��f˭�OHxr��~7<��x����C���[@�z��jT�ɮ�U�Zɇ��j	G��D�ZY��o�ѼM}z���j*����O����P���Y
��ѳ�|?��U�n���|� ��p��Zo��]2߮�w��5���'�EIV:X�!]��^*��jTI����J��!Q�q3����P�v�s�]��b����A�>�5ר��� '���x����t6x���Z�*���1�cȏ\m��m��UT"n��b(E۟C�U��~q`�������)�(QHBe�fү!��{w���]FVVAX���Nc�O��H:�Xͽz�&�