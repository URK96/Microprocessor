XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���x=�.�O��"p�*2�dʳ���f�L�	Fѻ�i�qTMЋ����hȊg{��u��~����t~�y�D���~M��X�csʗ���r�F�Bǟ��;�{�߆{
{M��wf%��������; �~���#ѷo�p�����W��^�6���R�$��LYi�֊X_��ȗ;1�}!�j"�K������pǍ��niD<G����q'�Rb�{�;���@'�_�`�_�D}�Q��;��1�4�Axe���7i=�`ԥbEџ>�c�J�d��:c|t�V
BRm��[^2"��Cc{�J����-�����GRX�ƾ��E@̭#wXR$�����?	�`d3������5L0��>c����W��d��d|@]b�^���Y>X�sɹ�a��y_.9g'����i:ϙl~6��"���^ل�>ڻ���zWM+u�� bxRd^>>�99�ޥT�X�;.jk�T��%�{�G��E=:�KFק�����T���|���<���UN���ze�-��=�A������9�[]v֏�pj�c�@kh#���Iг�q��y�4Ϸ�"����fU��Ϗyk�v���sn��z-��ߞ�W�[����ܲ�{V*422��"⮫���hWFz���!�)|��/7V�׃��6��������Һ��O��n]��FH�*oo�����]��@�� �?�t�oV��=�1�K6��/�#����&�i�O�z���X���Z~;�,�����EKS����`J7�h^b�� �ȵCXlxVHYEB    282d     8f0ҽ���A���$�*0Z�^����hφX8����[��tG��+���NЇ>�±$2i�*t�J�D��.ɳ!�}q�z'���<��S���]�Kj2Wܱ�w�8��KBD���E��2á�D����ӂ�b!��7.\����U�S�*lb�^�6X��S�}��*��4�G��hpKJv�����ZA#�~um �����8O(PJ��� �ɯ�:��ID���-Ơ�2�w�\5����1���ߠ���I�5�`�,�����w�SEf� <�����GP��`o¬�*�g��;�p���"�e��|۷.|;R�o5�>C�}4��N��|�7��GkI�&�G��}]�	�=&8~b��v��d�ԡl�����OP�S%՞t���l��H�5U��=�J���J�7�ѥ^�K�x=�P� � |HI	���5^�^wd��|���6��d��끈N��o4&K�,������T�H>A�*,UJ�<�nsB�Y���<8z����\|�B&��k�4C�2g97�,[���wL0LY�I&�xh���Q*iU�
�y���M�uR����A��\a��W!AH����4�3q��6�R�>���ҕ�4�.\���tY��噹2D�`4c�
�^����L��P\�AD�+޺�:|l��#����9�d�^Z��AR�ލ�����<���!X}mk��O�Tgj)t#�������"�ruĢ�.1!u���Ul�{���0�?/���@U 6�v	�b��>�vN!O�H|!�?Fg7�st��������L0/��T�%t�C�B	V���>nA�c=`������%�b�37�$#��|���&��5�fct��z�[$��qW,BfA�m�l� 9�@����L�̏�b~g�ί��cjZ�� �7��.��.|��^��g���.F������B���s�?����A*��WYŉj��t"1vx�!\��7��l(����[�]����o7J�?�7#��Y�q��/�Ai��P��b��~~��.B��~�Fr��{��.-�/9�į@�Ͷ�c���<��a���y�z��/��Y�C���^B��CQq}�d���)9����͖��-Bp���%������/�E���<k�T��Q�&}����:yoA��Gf� 0�_l�GU�Ƹ+��w1���E�j�)���XX�����]����c ZGg=��}@'�昉O�5�'5[��J.LN��~a�t?}�c��_L
	G 3j�S�{0���h�k�A�~����:Z��YES��V���W�Nk ��'ڛ��)�]�}���. R=���X������|h?H�A�H�S�an�/]b@ 1=	g���@+��W�������7N�������_\��9��*�T�7��XM���i�A\���eؖ�N1��B�0)����,ʖ�����"�.Ƨ��Q�	( �W����
�u����b	p4���=0�"�F#��tI'G�b�����(��#����̎�kjF��W�[��@�[[�b�pE�J��o��/W����'~�,�@Ɠ����c�o[���a�4��9�Rf�i�Ջ�[�M���X��%��=s���֋Δm�AT)◼���G�����-�=#���'Y��1��E'$~	��S���t�$c�3�O�Li	�ԭzq�z��e�ƺap��&)��Q�ǂ �MՃap����Fr4��ؖgi3+��������/t�'� ����h�h2�(R�>��)��R���"^p�^Xܾ�ҷ^� �}(�%��
$������qs��]S����e�K#!��N���R�sb�_T���qѝ�]xrB����[���*^'pM��T��0��.\��7�u�Y*�4��� �k��=P;$�oZ]����v�w��^��4��"C82��iSN�"Oי���<��J5C��)=�1�_��m��x��<t��,�=��h-`B5����y�b�'�N���j(�B�&�g�G�ƇaTh�����C�[�����ۣwUx8�^q>bjOT��ym>eZ�Z��f�\JC�Y�F����5�F�)�cҷ�M��õ�sA���q����1��S���rB��f������� �%ìK�[�ʭ�5i�I�U�r�b�����>.a?��I�2;d�C'��5�c� �3�'��|5a����nE|�&�M@7.�@7��wÆ!���Ug��du��p��5(Ē[����