XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P����S�% ��?�tA#�I�d�]�x>D^?��{Jr��Yf>�K��G��q���<��sx�4���� gj�p��\8$ߧ��'�:Z�������Pё�f���7z��^4B c�
�so�sȳ�tT|{l�Wl:�x����(Wg���(d�l�E��+#�j��b���d����1��I�P=�b8|��|G����+W�e|�c]Y=�
���A���A��9����0�2=�	��sS��Ix�LR��:����>���9�H*��ݲ�0N?��`�v1s�֝�1c��)�SH�\���	�\��� Z�;�$�ER�]}��ڏ�����Q$��%���!�lwQl9�;Q��?��	��-������0�`�l�e�?TMT����z�P)��7�w}��h�^���
j�ˠ����t\���h��Q�JS7N���JS���\���AVa#�O��:>rY��c����L��=�_�T�C�Χ�Q��G�Tq�'�1�S!�+�Rd� ����������adވ6���Q�d���9.á���i�:4�U�j���&�3t��E��M�rg�%�Dq�*4�ǃ�:XT�3��+$u:|��pNF1�u��B���#�W[s�'r��z @��'�kp�=�	o�6���v�eǾ�-vh��Uh%� ������%���j�>���&ݎO��\��!?�v�Ѽ��>ՉF#�&�*t+��~hߒ� WWHC<WW��XlxVHYEB    fa00    1960X����)�`p�t�����^��.��q�����C�G\)��&)&F��F�,�®ŉ+c�8x�'�yX��6�
���l1(-3��;�^E^"2����ik���T�,g�N��r�k������63��O�v�	L6���ƗF��L7%�=�� >�q�v�t>/�NU��Rҵ(�	�^�N�ƧK�/y�z��5�sgǾ��o1K��a����7=���N�ݯ����aW}��{�
=�Q �Hn��T�N����]��0ZS���-��`k��k�o�R��FcZ�2�߇s�v{�BE�Uzw�w���ǭ}POq���Rb���֡����C#Er5��'��MZk����¸%�-O��$ڔG�ed�����:��ǿ�V���J���q ��̀F�%�VP�ǟ�|�w�ChRD�������2��A#��$d�D�O#�{��ȨE?�7�o����S����铦��?���Aa���1ĊX��O�+��V�M|"��|Q'�f��֥V=P@�y����0:+s��U	�y.OC�������Gp���p�u
�k"�/�,`^i�/����?n�:d��~L{�8�O��։�w��X;�t�V������O+�x/��B)����G+Fgӻ�)������M)J�6xzg8�?�O��k�A����v`�D[����L����o�3��H�^����Zc�e��΍�_�얐�T�Fg����ڹ�MZe�x;n^�?����u�v��\��"�|sʱw�M���j�)	E˅%�7��L� �-����J�S�B�~I������H��ה�[�9��>�!�~	n�E��/��������,��E��2p��]X�W��.�ϫR��p��U���L��'%Y�h4�<�ߏK�l34�A,�eew��P�R[��`�+A���t$g�:6��'�1A'��0�6=)P<w�$r�>y�jS�,zT�2�\�{p�G�7����qG���R��Rb{|�aAG�������#�8"��n?>߆G,�e�h��	 �X��1�e5�#)��i\��K��W�~��#׿H���u9Vڥu_W��l[�S=�Vª<i��4^_���5z��5��H��V�K!o�?;G�F��)�hb�r���У��&�M��i�Ӈp��@�����al�)(�=��5m8�-���D^)�\���wIv"��R}��z�].�G���@{�^�o�NN��'�H6 ���|�.dm�Z�)p��d[��	`/���HJ�y`Rs ��Z4i��@�bmX��C�9�U�QJ�.�,T%���N+s�ʤ�IdC	�9US��/9��Y����A#�0?a,�'s
o�K �J�줕x+�ȝ�HR/�SDT�A����r�
a���X k"M;�!�4Z�������"�I��c릝���o�#��K��f|���~u�I�|�%�G3H-�yA�Uŏ��A,̀�:h6��a���!T��{�R8�F����q����l+���6e��o��e���C��2Moս�b)�m	�p
 yj����mf���X��x����/�A-��LLx�q�E����~�5N+�Ȑ��ˆ��C7���:�E�&��Z���[�k�~�C��v���>�8�����'���u�JU��s�*U���I�/���Z�R芢���t�*R���0�$QzEI	��LX��a�Ȟso�eՍ}g�(�#�2��٤��;�������|N���/ז� ��&��Kݗm6D����ی�K��]nV�sc.�������VB������ǅ�-�ZB�\������K�z�2�N��+f��ңy"=a�]`�������B�Oty*+�nL��c5!��E�@HI��x���c�C�����(P��8�'J$J0�ol��$����.���p� 8�wM$5�%�v�ÆK��*clAC�dv��י�&�����]�J�np��fZ���P<�f�b�R�G�i3��GJ�Ɠ����������b\���^d�{`����b=Z�3��٣|1Z�]y������Cf&�f�T�%����杴=%HV�Ӆ�,h��1�7�(�B�����]wϮ=�@��_4�J� �>���E%�����	��$��S����3"�hҲ�65r3�P�����{�b;�4t-����kTۅp1.�_jا-�.m#��ê�&$wi�z��$PC��P�BI��
���w�1�NM�K�.����}G�G�mm��ԉ��	mET�:�{���eX�~ �%�,�z��V/��GK����ی�<]J�gE���}�V|mf/��Aγq)�_RӶve!E��g�������y�d�Y�]]�O�|F�!_����8[�n��k��B�{0:�7�_",L8���6aX7�4��)��, 2�8�t!��vݳ6FRT�b>� �kV(�%�63���XlC�n/�Kb8�r�cHg���qX!+�Q����2�T��+�i#�l�Z^�X��jc�#�5��mi��>����.�&��96�����z������p5�����[��zM� �v��ت����?2<,���&�pq�1q��Q�e�ORVLam��+Z���ޠ��������c��&��R�4k��k��m�ǫH@�1p`#$`6#O�B8��Ť�I3%���_�V�35T����_�����.�����HmWT,f��I8b�{��������	E�������&u�|bO�&�!�t \&�L0�����+!�ej��4Y0�L��j��A���������5��9d�	A��j���^��Q���g&m}0�\ȢFD��g���&4G����y���x+\-J1����F�P�����h1�J��p]&ވh=��V�X�W���I��C6��
wef�>~�p����Y ,0J�iik����/�����J�D$�igC7����3�7��M����ĭ�|�f��j�n^��q�����!^�
�LJ	��
K�V����|�y�`�� T�!�z�
��@���\l��"5.Y ��W�Ρ�J��I`y.fI��d�Ì����-�|����H��qUi+�i�:���l���Y#���W��9l+sv*x
�.�r��>���m�����cI��D�Gq��L�lݣ>)�a��H�?���Z�O�G2�1t���HJצT�����o4t 5g������c��,����v^��~�u���������}gFUBC$1j�<����=��QP#�2*�2�������Q@�A+�k�d`�z�^Zۊ�1�{��HA�gu�^��Z��3��gH�o�?3����7��va�� �V�i�pg�/� ��ƒ�&%�e��r�/'�)�3�p�Ow
�HM�zN�� !�f^L�bń\_��.c��螁B��)Y1N����`���M;�`9�.�����Ĕ�pHXY(8�$�7~CЩ=n��æ��,f�
W.CO�p�s�J������K'�P���Fv�$E��(�?�.�O������N�?Tf\��]A�8S3�q��G�i�^QQ�2���ⳋ��?�� ��S}��zsX����U�He|�Ȩ ����jT�G���ܢ��ņ��A�Ka�s�U��Lշ ���h~*l�I���Y���L�j,�	>9� ����������/l��֤;������4�[L~A��;d|sXÚ啺O>�`��5PX��oh|�Iq�6��\��bOr�1B�"�E����V�����iPT^�������=[�b�#�U}���Ej�9���E8�س2�c��E�kW�P�|��w�������8L8��g�w�ֈ�/AB����� 8֮4�j�'ͿȰ�@L�����	��.E�k�6
���gy�k�AOi�8�W�1�d�#��G<TK>�;�n���U:kcG���*�̐g����<�I�$u��.v�t�p�44��/�;W��`�������dCa�سͻ��~��O��3d���j�
G�}�`��l{�?^�����������6hWO�>t�U��g+�Md��3&}x/�w�x
���{�t6��W� ��rL��f���_���U��e&�Z����u�5R:��YT���M��:p�0ȯ`��L��;��ߍ�@�t�T{���c�Bjvņ�"wP3���'�R��c��K�F�Щ�����b��6f��_ռ�)�KE�AmR��Q��f��td�g"����FPp �Ϙ�Awԃ��m�vN�o=�{yU�ф���A[�C�c�,�`ǀ�Y��5���n��O���Sp��%ӓ�ձ�yױաi��Mt�U5��s�\������ڽڙ�.���쀮bf�� $�x>��/*����4f���x'�>j�R�����sd�P���ǅ.�����������_�ސ�%.aq���U�QGA⹘�WrB@��������x �e"���� ����'"��@|䶆�z�����iE,h24}�RC��?�|j��z#fټ5N*W���g�x�ћQ���$N���Q����9�My*q��k,.}ym���^n8���z"soj��U�k~��Cn�j��]$�Jx�n�]f��zE1x���\m1��N�"��)�ZA*ѷ�����ZYP=X�y���L>W�ti:��{�7I^C����2��ڃ��qr���iM?Pa��8���3Fȵ�mK`�5���\�����},ѯ��)����=!@�ne�rD��"�����PЬ'K�($�1I;F�n9�t֊e�Km[�y�����m�����`R�z�R(K�]
DXt��.�LIc�`H>�+V��E�����B�������v+��Cz�C�b?s�߱���ix�X55�U�L9�6���-]�l^';M?�u+%cr}�\��|��/�U 5{P�_а����}4��z[I"���'�zb:��K%O)3hS�S&��+�x'�_�z�ª�\����(u��i^ç�9[�1B-��X�,F��]�5ՠ���W��x� �u���r����s��5�ɾX���O���c���D�4.!���n]¶��q�m%���,�Q��Li����>p�`�p%bJ_���+�����C��-߼Y���j����wU7�T�xG(��6f2x�.d���5j���S������dS+:D)��O�Kt�v��D�s+ދA�t���Z2X���RYr��u�;У3	�`� ĥ>�k��턺����:�iݒξ���&(pVj��~ꅩ:��4sy@�yY����p �MP*fu�c�ѻ�J��-��~�Zx�9.Raݔ�{�,=(�
/������&{Ɋ�"tx��%3rk��xM�b��0��118�����|�b�35��$Lp^��7J���25�no��9n�:[Bq#�ߗ�e�z��\�4a���2�	�䚒�M:s�B�(��Ex�q�*��,Pm�ϣX��*�Z�z2�0%�}MݽHo�X8�n���:L�~��Up/���8,X�[���A�d (�u�LxV�������vEӓ�(�|'
������vD�S�W*�N���f����sδV�������Ę!�T��嵕<:�F�F@h�9g+��6ӕ�*��4�/��3��!����u���{eRےB� 4���m�@b��+�Ko��H�y�$�D^n�3ǋ�@�k+t�����t�L
i>���L��I1��.�D�ml1T�@�c��JS8{������O�.<f��+ͨ�����@�nl}�B+e��9��u6��w��nt�#K(�tH�XI���=���>z�Hj���s@�!����xP�Sh��f� ��u��y�ƨ�\]�f;ĭ5�Ii�M�Ev-�h�-�MR ���%��*�0��$y�5�/KR��C��3���ܴD_OPl��8��"<C/���儕)( ������|�$ 57e�d5��Uŧb�w��Q�0n��� EJ/�(�4v,p���h�9X�d��uSx��6,)ۥ��ȟ��l��;� /�t���v���U)��mS���0D��D�fV�����#�&�U��d3����%Žy����+z�}��
Jh��Y!�>|m,��-�-ۢ(ˠ9H��g�M�В��(���|`|72�lX�i�;=�fp����+i.����N-���>�q�*L6�r`�o��f�.�q74
�@L݂���7�H�Z&�'�eɘ|�p���/�k���x��=�k�m}$�(y�-�j!,6?��9*�O����\o̾����� qp܃�5en�����������5������"�������|�$X�PQ&7�c	I��Hb̟���>s���L5����05s�R,H�V�b������łwۜ����5�F3����m�	m��`[�=ʶD˰�Q�= �qx~��x��(i��#��S�����b��c�Ә~`'��XlxVHYEB    fa00    15b0�P�[��%렋D����cAe���pb10�-���|f_y��^#s�_���j큠�J�6J���s�S�K{X)c��!F������ܟ�_����Ɗ(.��_cG?���e�R���x�O6g�P
�u57�фv;.�ʰ~	|݅�*OtQccc����z-?r�Ό��elK���*ࢼ�I4%h �����	�Ȯ�� ϴ�9GĞD��[�4��~��5����M:h@mL��J� ����t��`�{W�񭹍�e]߾^U����0h���'���qy��LA���T!��ԃK�xڢt�H�޹نS|xj+�@��	�<��8���`����f�g\�r>d���=��2/��&R_�W�|Nut�#"aF�}~��!���_[��7<�Z3C�y�j�$qd��l��jTr�=�ͦpv�A3�˄8߅q��cv*��HN2�I>S�E�L�/�ޢ���Qgh��ui'. ��R��m�&����(��k8��hG@9����Q��@��]���L��`�s�{N�G�F`X��0�R�)��	'}F��X���'2C܆��&�$}i����8�S$L�n	��b�M��EX���Ɨ1b!�a�L��+�i�rI�~P_*�\9_$�h�ⸯL@��_�A�t�\35|�ݹ�k!s4�|I(���^�;#2�OL�=8>P[�����I��F�+�}b&B�|$x��c��$��vz�k�����(��@D]53��":�2�wPe��<���|������^�:�~�y��¸-G��c4[d�kVr(3�:����sF�e������\��9训x����a���1br-+�ы��K	��ؚ�K��bR�G_}c�P�	s�?��{V����v�����/��$��1�X�}JQ�4w�iuE�c�4����'e���o���I��?(НC��u�D$l���ӡA`�0� ŗr�HJ,\$��2[uێ�s�q�o9�� ��k�OE��B�G��Q3� %��g ����tu�$�:X~�68'd(�HC1c_8#����6��6�hŎ�Z#
��Y����g���9}�i>Z����Ll \�7!�������9�{P�)U^�B2�ҿ���Bf����D+�E&�8��+\�.ɞ=ʅ�N�Ŝ�MH��}]�oˬ�����=ۅ�6��/��������@����+�XM��/8Z���HT�)��x��̔*��A�����UϤ�g����
� ����Bm2D�!zR>����"��1<K�N��̉C<�n�^�Lu��W'}����ʲ� 9(o9��~� 
��c��Â����
Q���H��dC;�}���Ty;:4n���������b�|�}�G����.�Pn�~�\Vr=b|{v.z�"B5<���j��Bc͗����՝�g��Un��LDN��봡كZD|,ї��5?�C��z��a� ������0[�6��\~�/�����^��>���\g����_r�.���?���!�����Wt���\�l�Ϣ?�f���C;����Z� �|�'S-����N�t��B��3R�����>�]NTгصd��Y�O/�E�rx�^>�����[����2�6����A|9C>Q�=��:�2C�.���b>�mY�m#�}��ڄv[�ktn��k,�ݣ#��)qp�!�a��̿X�D{����W�c��4oyi�/h8<�l'߂�j{�n�7���+�%o�6&^����Kv�S�����
�;��V@\�c�n��$�0�Q��n>���|\����R;nqd^6.$�#%��;=�`
�z�|�R��y�ߐO�(T�ˬ#�p;¬���ӜN%m(�?�9�=���0�+�l�Q���x#�]Ej�t���|͉���U\��^"ՍYBG���Z+�����(�3�`!.�"�'��Qw#�B�υ0���n[�!@;��#o��IQ+)Jғα �Pk���J{BH��x1��8��򆏺j�7"��Xm�c�(y��*F;��7�������?���R�H8Y�J`��%ގNf���U� ~XW��Qg�(Kn��Tw��E0�qIF9�|�!$t�/-���!� ^yaz)�"�JK$�7x=@ܿ����N:��XH܃1�wP�vo V��Ѷ�yO{����f����N���5e�c���t�*sq��hh%����t%�L�z�]�<��W����ca?0��7���l����2EҲ�稍�>W�0��ӟ ���`�F�VnM��rn�	j�p���U�fg
�K{�l^�����r�ڽ����n��*4{���۷�iP:^��.��D�!V��ctF���C�t�La���ѺFe:zF{m��>�+�W�k�W��V[�
:�t����7r{��
�� �'4�?��2��Χ���%��	~��eˁ�R��$]&S%i���9��鞙�Ő�	t>G%�������b��(�rPJ�u����B���(�d0o[?��c�ю����nv 7������`��%|�]g ��Ҩ���"�H�ebVI&(�:LԜ!h�h,{R��l�3�Q��m���r �z(2��V�1Fٺ]�@��v�4Ѹ�@5�&x��v8�e�ԖMjOO��K}_��7�����m�c�a���ۂc��zњ�� ;��2,ģ�f��C/.����]w#k���cK<d"��	F(jC9B"#�S�[��D9��bR�����v��‡���lӃ��R���<���?�2�>��|��X�"���cb�4z��fMUR,�Ղ�H���z<����u�|[���^����9k�����"��O��m�uE����?2�VUY�!�w&�de?Tn�+�៸��额��&�`�vJ�q��Pڋ�	�8��Q�b�������+N��@�5e<)���w�Lu'����%2'[�[$�����k�ȼp�Iz	QxUuؒX�Oo�"ӊ��9 ����7 !#�e��ޠ��� �D�X֯Ȑ�<>���翱�G4�H����5������������<CW��$��h�X�s���'�ζ`e���iY�3E������'�;�����$�\��r�&���A<�r���?Fma���zQ�4E�7�{�i�( ��r�CpW�>{�uZsM2E���-lHDU�u��
(�Tb�[�+!N�["���MX�)�Q[�"�l��+���hf�6���T[˱�eҮ)5i#;�]�����Pr&��l�R��S%�Ƙ���`,s�-^��`8W۸���d�bp���Q2�8�钕D�Xjܨ]�=����W��}D�WH����1~1sS�p0�����"��� ��m؃4ϳ�������F'�<�����6l�˘�=  �h2� �V#��`�~ߌ.��2 աb��/�&r[�v��6�jmmai}]�jGR�,$��t�4$r+�W��@8 f�0�ٳ[nA�RbQE^1]�j*��@�h޷#�xƻҫ7x���5Z�K0��҂��<�i��SUTEp�������d�{���_��Y8�\M�K����z̰��W(<���uu4��|��Y� #e��Y�Ɔ�����c�[W�^RO���~���d�iK�;*�{��[�s�CY�R �'�(�|�[�f���xh�G �M����a���A7�@� ei[����R�s1�TsGtS )�4�$��gJ���m+ m�G�1���ro���@L�a��$p���y�$� ��E}����`}1��l�^��r�1a�Uz:?KC�����Fod�/x�BK�ÝC�K㝇������04��Όo�<� �"Àr�Y���_t��j���8׵��B�p���Yl'�BƁ��A&��o� ���N
�.(�&x���S�>p��:�-� ��ٝ	26����/�I�����<�H��u��b��w9���E��t���#b���):\5�������ߠ!�����r �	��{�E6�ja�o��CD�g�Ax�3eh�-�9CA�5��c(̯��>/���4��j2X���baj殩����Ţ�;�~��[�r~�n I��v��ZT2{�Wƍ$�� �-�I��3��/�	i16-�fv�������J�eO�'*}���l�~pf���(�"LЭ�z����Pn��b���?lb�	 ��M����I�}R�/N�ix�9��5��b��k\�u�Ԥ&�TQl4�OF�̛�lpԒ̀�72�<�3+p Uzv�7�C��C���锧��Cx�@�IC�أb��V\+d\��(-�`E */��� A59�51���Q���y�ŷq�k�)�.Pn�ع�0_K8 �������A��}_��p.��2>j�Vad���2i���6dN��?	Ta����Vk�T<z��z����g#/�s�# ����2��N8�!ޣ��ؾ��S�����v��77�9B=c�߃?�e��)Rv�蔎����9�����e��v۔k�å깭g�1��S����=Nd�M��{Э�u�[ެe��ǰ)ߣ�����-�t��8�ғ!M ��dU�����:�x���X�"m�x	\������J���۰�̮��鰔IX��9U^u�g�l��w�v$��E�4���aˆ���G%'���<� Xe/S�u Ծ�^�iX���^?����bU�0zi��,�߆���9�ބ���]�+�U����?��R�
�����(ER�[�8A7�u��E��Nvk��]4��4�Ir>���T(��E%M��0n��U^::���o◻rL ����('-��U���	|g_��ܮ-剺�w��qck�r�a3�q�ҙ})'Ȋ�ɞ�XN`}A��g��b<>��m���h��
I�[I8K��5|#���S,��.���e�J.1��趮N*����Գ��f�b�ټ��aۙ�B���dAưA�Y����7���ú��	{��)d�u�aǦU:�C���p'59�F��p%���N��.�e��o�E@︚V����m�)�)�-��YI���m�O`S���9{@�����v��6m���"�*�x��������Y��E��P�.��������.J)]��^<~ �|:��O�jZ4�mPP!��Y��
�6�tWl%_
��y9@�ì���i W��qbDRb����w�&Tԑ*w�C��� �g�4 ��cЙG�i	�Kp�'�' �m��-���V��^q�Ud%�>=W��a�xR��x����}��{��QV��spz�].�2���}4�X�=�����۳f;{m�i�.)B�LG�~G�ĸ���#�l�@w�h"�,����]�tg�f�^����J_��J�CA����a���T�\4SҢo}i�Fi�	Q)f�C���:)�L*���,����mx�$XlxVHYEB    fa00    1600]�w�I��7)9*�Q��JH�Gx\<�(�O�Ắ=�|���u2E�N(��:��U������~n� D��Q!���qнQ���S6���J=Ak:TP5�Û'�Gұ�
%��0~��{\�2�~��m�]�J��M� D�e�a#�t�� �݋+������c��u���7�E��d�����8�i�)�m�E辫�>��ְ.�����q���c���h�H�ˬ'��;�b9)2�m��:t�Ҝ��8���DlN��^��.Q fu)ʘ-��j��0���ΰ艏��i-��럁�1�9&������:�(�+��0��y���%�Bˁ�h	��O���Krd��;�G��֩���e��];����Y��7pڢ�!���~��ӣ-�/�)��/W!o,_˔�Z-u��D��&k?�Ye��E>���q�;KR@��ȳ�k�l��zu�`��7�H6��c!��C����)��ދ�+�,��㼊GV_?R��^��y
~�U�#�{�_�*�ia���i���<�%tHL�cr�@Aj@���ڬ8u�)��"���4�
	ݠ���ö�"��-}6B�&H%�J���Q=R=6�n�kTg+�?NG7@�ۯZ�{�ei�������r����8���irҁ�F����ڽڇ�M�a�(�	����Wӌ�}�r{��_�܋3 d������y�Xx(f���t�|k�8�郎&0zr������F%�1 �
SA�j,! �-�3_RAԵym[쁝�j9���2.��<�3?��D�	�^ח���(��9���Ti���re������*���ԣ�@i4k�'�E=x��P
4�*U4���.r4X��h�h��ǘr��P?ď�׌hV��*Qz���+MlN�4�9��^���䋱	n�D�]$��}EH�]���H���;�0j���xu�[��Oȗ�v�T�>�{�P�� ����dQU���
wS�i�K�~�H�+��j�޵cJAX�]����
YE��� �m�4F*�`���>^�S�+��K��M�l����*;���2U��K@G��krB��r{<$~@��5�9�W���ޔ�O�(�B+A�i���}����f���4����6�0�V*�9#E��_�3��m�\y.�I{��8iv'�i�ji�T���Q7b�ˤ�Y�s0/w�G�!.�gڋ�.��y$�`��#��m'&��Y��D�ӽ�S����m�ǩ 8`оj`��H��X��2��YVt^�l�������{�����
n�\�ؕ�0��d��FY������7�8 x5fO&�3��#ӗ�s�1�̉�1�a,��2�ub���%Đ�0�z�I�U%p1:����`[��{H��Uwt���2�l0�a0���ֳ�X����"�$��\'yj#��$X�He�z���lJ�1��m�;q��`�+��x���
��4pY,�SP �;]�}���:�+~g��)�Y[r�i�Jr-1y?����1����9q5���i,�{Aa���5{#���!�t���O��9��V!���T>��n�cz_��G�#���d�yM��䡎_%�?a�7�u�* �$	(������,��WҮ<��s���P��nө:	l�B�s9���/��eK@;�m��:L�Sy���o�|���6�yN�-%�mv�L�e2�-D1�Eg0ns}��qP�/[��N�p��j�<���Q6���TR_a}w)��8�Of�*-��X�ߍV{��Y�z��Q�~_�-g�=р��c�4���#���5�}*Po��v�L�eJW��>�c�f��K>Gq[�YP��z)(��ih���(��6���Ҿ=���K0{KH����\�+��Ir�3���~;�,�r���,vW��H�pof>)rB���m;	9�|��ϧ���Y��n���35"Ҿ_��֣���2ĵ7Th��Ǿ�*��#����u@�f�N�F����h�l0��D���������Y�����0��o�����EF��n���Q�ߵ���=���n�&��uR|�	��ii���+S�ՅA�
��q\|9��K���Qًcg���T�t���e���gI7���8)"�c"�ʹ[��_�h� �w¡��s�����U�?ܖr�y�'�{ ��I��?U}�h3Q�|y�HJK��P�?܉�\���ᄥ ]odݎ�*����Q�]��j�����=�_�.B���9_y�ZF�w-���Gb@�^D�w]m�챰´KyY�9�(��D�)ǩ��̨�d(�[�� F����9x�C"��:B�V��QGk�{ri��,#L�\�cO`��aH����zW#i�� bpZb����H:3V�{�so{Q{�	^" SL�'i�WuJ���u�N2����d�0���O�&!�9x��O4sA�e񽋚B���W���|��I���	B�$�$�@��`� �t.�M �6^�_���(�߆��D.r��)S���[�c�'��'�S�b�|h'��1pLn�ų���+�Z����	q{AԖ?�&ٛ��6��	�&VҤܜ�i�@�j1:��*�7�<0��w?Ƹ���.�a�m(זTT�VÖ�
��2�e<���^���ݖ�I�s� a�)f�����9g�e8���4y���:z��A0���I� IH/%���CT��6�Ie%��q
��ACT	������;R\�I��K�\�6��nŭ� ļ�Dh�؏"Y��&�@�.8 �CŮm��K8Vܑ�$�Y��DÙj�J!�f{�$W��}���s�j�`��Y�O���V�w������2�p��n/C~BA���>��K��������KLd��(�Ē'�����r�J	F��A�N��_����L�����6t����}�k��kQ�6̓XH�8�<6u��i������l,�h_�ׁP`�� �?���iꬱ�pH5�,��G�����@��wͧ�Pw����+nB~K�0
|-�gg���Y�-��)|)yIv�����Q7��mr�8��.:��DxΚ��_G_� �HW���;�י���oА )�Q��0yT2a
��OBj�u�i����K[u��I���s=���qz�㴂ژ���B%iʱ�&�Ț��Q��~�H_��vn(#����Zb��Dk�t���R'ceֿg�W,M��߮��`��	,-n���b��K�q��&e��hYa��!�O���,�:X*�h��<LDvth=0�˴��y����j�K��������v�vnzk��0S�j�A�m���r��h@Sth.��J��m��r�E8�'+?q��c)����:����2��?�_E?�>�Ae�IU�j�b� E�-�#���L���H[8Ԍm����1}c���!C�+G0U��?���H���@�CI��x�ѱ��$��K�T�zP�y���Q5�2��j�C�a9�%�;F))� }��'5o$��U������P�K\�U|�Y�lޭ�dR�z1�;≲����^M>�<��\o|T�2��!��Nv�&�ab�����eᱛ������ =�����q	����t�2�1EW���Q|ΔL��ZҨ�^�¢�o3�2���L��~�k�e�#O�!v���ԋ�1`����S����������2�<m�o���!�T��QLD�H�=�-�]��
:�@h���
�8vm�O�x�b����&��ߩkM��{��}?�,��b�b��3'_���!$z������7"/,�����rǎ��Ӟ;e�
N�u��tr�C�l�S�h85���)��� ���)ÊMn�e���!��J�0��>�ƃ�b�'N����MO��S�c!`uk��G��1וwC�u��k���"�r��l&�w<��E�� ����sk�B�
��A�Ė�P^Ȇ��p�rkÊ��S�f��e��0��l3�߶6�^/��l���C���cH���3�x��$Z�K�����0��Gs(�,F�?��۞�;�m��/~����	2[�������7�H��kw������D�ԡqD*}4�H�`�r�ڧ_� l�U=��,����xf�fޙbJ�t�$�eu�$O���o�Z���g��v��Q��3��<o̪���e,���I~�6��c����&Y��S����FA����Q�PSɢ��y��#�]b��VP=m]����z�n`��%=�[m<!�4��2}��!e��6�*��_�;�0�,��N��X�^]�Ҫ��:�Tk6��RNM�I1�|�7�S�&��+9O��R7)P������e$B�Z8�fS�㔤�NЙ�^�/}�@���lYʞ�!�\/�p��,���>H!t�O3�چp=�]ts4�����s	i�M|:�v�>d3��H��.��'����y���kLpے��$%]S��
)�����&�l̬���'�(�~Uq�b�u�a�!�;&a�bm�ɒpau*�9N�g�3C�I���17�M�x�|^n�q��F����1��x�H2���[eϹL���?�Өݡ�D�9��ݖ:v�nն��wy
�h��^��P���0�Ȩ�xf��y�T���R��vY-=�}#j���J��}��BP�u`-!v�D�[� �����ǹT�R���N0����Em��/ @*"F��U�<��'�ـ�ڝ�_�M�ͷ�9jT�9>��8��r�Nl��y�}e���X'�|��Q�~	�8�I����(?�H��a�5�W5ȀC�0�}�ƟK�ĵBf�_���ܟ�R�Ⱦ=�o�E���� g�fL"
�E�ξm��p?+�*�Hg���nz�4��ڙc�|��'A���w*�3ܽ�*����Ҁ?��2iu�첽_�f��ô�,uPgn(��
����ޢӕ9��-vu¼���D!�s���*98���c�����zhmuR��y@�3�۽��b�����>�-����~uAB��@���9��O�&c��OU����:��ᷓQ=@�Q�-+����Tc��Υz�k���\+rǡTX�D��	�s��WW]�7M�,k��]o�&j(rӶ��ʾSu��ثg��$��/�,��)�� �~A����������#�rj6����8A�	:���c����si��8����^�XN���A~��һ����ϗ���$�ߏ<Tm�����[j�U������Ñ��d��Pr��Dl���0�Qwb��J�� ���=Z2�A@-E�ݺ�#B.������ڐ� )}�I��w��� W�_*����z$ݫ��#�z�����H|�XQ��D���ȯ����xCl�LKZ8ҷ�th$�,��ٝ1�����x���{mN�(�Q��!�@�ߦ<u�"7㏒h3��B��3+i���>��H�ލ�Cb�0���b��:�P;�,��6�霛�Қ��Ca�;�v"�X��u��i�R��Cz�y�5]�_��%��˔PΏ^lԲ+�y���l6wr�����#ή����z/��$`:Y4��������)�|;{�/ր!U!~)��V�`�ƍ�ڋ�������:ËyꤵXlxVHYEB    fa00    1630&<��d4�k��﫚P��Ȋ�!D6T��f۞}/a����?ͩS����m�ԟz�۹O�	*E�Q\&翀��']w4���w��Ue��v<����nEhfy���iZ'�{���f*���L@f[8�VR����:�!���L��]�v�b���lۀ�����Pf-�poڞ�t!/�#n]��Vl�,�`��-N����R�_��pG\��3���H��w%H�mNd�9'h��X��F6�+���vO�P&d$���>��;���>�B�/�S�����7�sR3�mC�O�a�����ݹ罩�6���ȧR���AΦ�� W���I���]r	-O.m>���qڅS�8��V�7�&��=� ^�IP�x�J�uR�`�]G��t0;�ml$�z4���� W�����D�dJ�O.>T�s&i��O�O�`W�P������(������P9�\Rk��+�ܐ��BwT
��]Pe.�����7�����:s�	5I��BV����ـ�*����hb$��M|��:���X�/�Dl�L?��㽊��Uu�;��b���R�f4\�aKݵo��v4t���s&m`(&|�BB|�9����5��6u�n5�7V�ɟ���Z�&��Z��l�
y!�s��N��[�ݛb��O�S��.e͒�K��U����<�͆�v~�D��K��k�Q��B��)g D�a
��{����>�'<3�G�>��?9�Z���s3�{(9Ґ�ST�N�m��[�j���5�3���@FA�H'*+���h�K�u���iH,�����%�N���,�����d���K0π^^������V�3��%- �_S�
���*J�Ů�pKJa����4ċ,p����-Rs|f^o��� j b��j�Im5l�H%����fz���
�7w�'|Q���Cz��F5f��:�Of�V�N3�k�'�9)�GJ ���Q�V���ݠgsG�*p��DyE��z�{��G
(��cݳ�y�s0�~ֻq��eV��*��Z�n �OV�q����<�q���d풔��R�l��.ׄ}g������hO�2y����:���u���O������� Ns�+��6�;<�z�^�A�'ɴ.����0I�����Im���VzK�)cۇ/��[79y�f4'Q"�Iݩ��KӸ��d?��8c#|.��d�Q,�rF�SA|,FʌX~��n30�f_�������?�����OQvC4�M�Vrڣ&�S�3��/��HF�n��#��b�j�$�D{��k����l���0�AK=3�6O*(O�Ō�Q��q��b�\�����U��W�o	�T�����!�V�y�g��v�Om�x_i��AT �a�ρ�w�e6c��s�����c�+����Wou�J�,����Sm�I�%4�}��M#�i��٢r���XEC'L[`:�<����-} ��up�H��e�����i��QmssS?�EA�}�
�l�����"���c%N�Q�A�/p��P�b�Z"�!��A�I##����v��nIܒ�CkS+p��կ���b��6����zW��8s��b�E�?:�ԅr�I<K��ká��ǈY��`j��u{��Eƴ�a�q�D+�J��$rɞ0�}�![@��Z���#&�2�m<JH��▄��JQm���������!���M��(�.2.���(7a]��_��z�(N�LJ�Z�{%���q-O�%���;�RY?wc'�O-4��[s��zֺ�I�������^�U���6׭��� R�M����f�Yl���I9�!�Y�r�`�~xT��[7˿��AC�i�������hLd5 6#Nyvὕ�T�J/`���%�o��.�bl�씬�q�C,��Z�B�+5�F[���P��ctL�^d*2��'��#U��k�ɶtF��t^LP4?���Z�
�l�M�Ol|Z���*h�W��3�0|�֍F��	���:*� Zɇ��F�@g\C�$��](�&G%�ɐ<4�֦�;۰\�v��z0p�z~��]�l�	���e?J(����Y��:uvm4��-�u�P���)'ܟ�3��`���h�D�'݀ d�^�\�`�2��S����d����C�BnB���]<
��.�q)��Ӽ!��?�q�(m�5H�kl�X��ёK��{�g�khL��D�����[擀r^k]_��ռ�o�9-�'H���;��w�#��!fK�u|�<�Z	�Aj2j�D���<cg�-��������73�����i����Kl_k�6�8IH��<v�q�_*��YpggT���4Th7Wq����������w������U/^
�4o`�y�솬U6�de�yAkUdba��}X��x�F���l�'�"�H�I���ڿa��{�j�(��K]+�0�&���8�
} ��UY��|5D�!��ގ�BsxT+�dA�/�� 2a��JD��޺ |�Ķ��9ܺz�Rtjޱ��{cѻ���
b���O�O�' �Tx&w�Ā�dE��Q]�N�! x���:Y�rLnO#�c���tCa��	B�������О?�9�h{<�K?G��T��΃�Ah�PG�Q�\�
|�e.}�0������Ɗ��/轒A�����$2})L*B��f~$�X���*�O����3�Ԟ�#
����t������x�!�;Qa���?�u*4�W`��ƭ�6�1��G%^�+]j�ר�t~�k�GAbk���ǂ�{$�җ��/�"va���Ԩi�|�YI9�H�Z���S4�-�I����S�u㌙�BoW���:�� �N�����ɝwV��\!
$��;��g��b��{v�(��nn�Z��?��n�����$�D�/t��Y�)?��F[�Z˷�{k�w��P7-C��1Bci�D��H��M$T�Sn')6ݶ^�	5�G�@p.ܧ�**p��*Ǉ_^oG�OA��L�	4*?�R��[���A'�S{Y(���Q?���M�V�{�;� �xe^^gO�DQ�2�#g	N�=����=n�:������'���/�FH@��^�]��Q�/��}��@�城�o���>i���j�^{�p��V���ޘ�染��{q/�:�;p���S�utAo��{�=m�g��1]�,%�(�HBy'v���lx}��q�\��-N%V+NI�����^e��mUe�j��[:Η�o4��5Yr�F��-m���2�Y$zQqĔ��
�'$}�;p�K��θp��q�R�%m�6��ozaU���/�/�Oʫp��v�H���;����Z�2�%g�!�رǥ��'Tc�rǟ!p��0����31����% R�Q�7��xdҩ�|�OE?�'��˓�V�Ob��bG�7�IJ�K�4Z��WB�9����4��m�xץ	���Q�В1`t��ѾfW+'0Eф�/�����ڜ�
����}E�;�!��e�[f��V{��|�(LI��
�ӭ�}`�Ѫ8e������k�����Q���?��g6M9R��#F��Ͳ4���ƾ�H�xg`K���Oω�7�W�=zU����=��@��B�K쩌1X���l��^e..�s�Љo��>���{���dLO�TO|:�~�5G�����M`\ۜ�X*\\ߗ�5p��.��Ct�Ͻ�OKE?���7A]7�((ʒ�z�0�%;ȗ=�5�3S��Oh$�[?�J��f�=�X��=(g�.���Ow*ѽO�z �M{�L�W���J8f�l�}u=f �c�qU�)qk�c4�^�p1$�HXx�"J��D.��$���V EF2n��rQ��Vt���v�/����Z�h侉����:ćI$�����xv��bE���n�Ԗ� ��_�7�i	'S7v���y������dy~�轥�Ɛ8���"q��v;37Q�u�LS5�
������F��l�%���x��|��z���H���"W�ߝ��ˉ:�y����S���p٬	o�/�sW�`]D�ղ	<2��ʃ�u�<D>l:������^V٘�>�a�u�/�l�
��z�6�.��e��8���=	=΋
��o�	�0�?��x���!�i�\m�V)�9V�x�R��J�^,^���p8e���J�|o�	P��(�JX.�ߚ��!��+H�/Z��OAoo��U6����� ��J�?@yD�#l*��6T�ؾ��Z�>�RH!��H�[�d��R��g�od�Q�@���S��f��H�U	�E�dW��G����U!n.`9�6��e������2���)
W�&?�)�����tPoRoa�O�"��tT�>���HX��s�  ��=��/��p�9����>)���53@���EF��f�@�S�ݬ�&�0�r�W*��1���������[(ȩ�^$���O��)��h��T">�3�-�	iE��B��a�%[*y�鹄A$�<� ����0?�N�fhxv]������6�5>�|�Dun��D��[�
�� �Eb���3�4�����0շ�{�����/�w6.�5�/�15���
�2o���g��z���.?=v��U'���.*���mn3����i�f��
Y ��USt|&�/ע�J"�Y����\��C�*�W��b��sّ�3X�C&仔��xw?Q����s!�|�W���ySlO3�~z�O�(|xB^�	�T�.��9yņ؝�� z��`oRɣ��y�u���A�)'�ҙaV��U���ڍa@}^BG���f(#j[�d�Yu�38�6�5�͗	�Q������A�
|J�&ۂ<D͋7�h�ӈh-A����0*!ؒ'yj`��0���_���˶�Gߡ��!#�{ RX���mѫ�4�L��-�}͎C��}��9��5xf����ۤ?H�Dא�@�e�<�涗2��~�t�X�����Ħ�-t�*����%|����_)�?�̜zx��ZA�u�	����񃩖��˘�(w��PZW���i�P!v)X Z�
���?��t�)$UM���C�ƹ:�F�y�+e���F
U3�\�$P����q7�������&� Xs�l~�9�"X~�7uٛf��cz��E�����g�1<���zr?����Ws/vad��̣y��YV���OOߴH�-��H	�P6V�xq��)�1MY��w7�p����L�W�1�iX��C�Z�U �rF2ܱ��^�\��XL`٭Jԏ��a|�S�$Ĕ}�9�����:���r+�� �Ρ�c(������,Xl���N"9q˃(B&��%5��'����(W�M�3��Nnl���Q���7.|��1�
m��Tʪ���0�/��'�?5��d� 0��} �q6�Z�C2\Ã��Oݘ�ʻR2��Yҿ$�K�=���G�T�4O͐ۼ���E���F�q��+XI?�p8���sK�ƅ���b%���Y]�D��<c��H��F�������^:Lp�\��{)ɴf�9�G��yX,���xI���8M*�2Q��	J!D�����<;�
/+�v���"aA�������T�׭k�!���~bs����v����?d�%)��C��b�T��L������/WAZ��	T�i5r��dXlxVHYEB    fa00    1620�X�hWp� 0���a�]B�VS�v���a��)�:浅��F0�������UJ|��L������:|����%�0)fS=���c`wN�����L�'% ˏִ9��
�jx~ѫ
Y��^�q� ���hW���ዱ̂�터�Y0�6��<�I���]z�H$Ꭵf�,t:U���E�N�-"�^�$�I󍋱�J�Mz�$I�� ?� '���qS�Vg�*,9�~���唐&��e��9`�2SF�B!E��Pp��0��n;�
9D.ɛ'��oR4�C�əU�k�P�P��t�XF���Ы���D�s8a۹��J��P����E�p����~	�A�Y9�p�S����o��u���|���8�n��ZZx�u�av����Z�Ő�|��F�z8Hw�X��-q�5 "�M@VS2͜���X�\��(@�ׯ�`��!'�&X��'nZ���h��$z�D�6cy�SI�\��Z�g	���|K<l��F�n�\��w��B�8�!�T���ϕ�-����@A�J�:�0�Tlf�X��Ȁ��guWB�L��.�S+��$�bܙk�G���C�ͭ��+Jz±�2u�PFJ�����
`l���Qj�`~�<X���p댔ya��`��4�Ч���U������^���F���[*�Ȓ�<t�=��q�$wݰkQ�`��w�o�6�3�1Jo��`Y,mQߜ��o4�c�>k��.!�i	~�pm�@���-��ÝP���4N8�ucl��?��������"δM8;$9��jHִ�.S��8�Y�@����v�k<����O�9���ԓOo8T$�ia].���l��D�w�~�͸c�<VE�pxI� 15�&ZV���\�
����%�TҮ9��c5L�EO]Bx1i9�1��m����mAl^��!ʖ��>�m�K�	of���8�q�a��~���{}ߖ`�#B�ur�r��n�����$1�yв��d�t�L��Y�،�(���)�}h�Pv�˘uHλ�%�^ X9���3D_��Z�'fm��&R��SŪ�v��� �! o3P�,�j��6�j��U�7�l��?m��q����*w�c�X&@�������c7?]pM5|��v���p,;�!j�I��I+�7��h��W������m�����4j��Tf߃���{��{�֏f��ep�m)bζ�u GxYx�[`��JM�2+bn-��.�?@Yd�tѰ�|�苫�A�r5��*)��!�ئB����%{FWZc�ܜX��)Jqe/�!D!���w���� s�T&k
�f��J���A�r�H�O��t�(�	�i���u���{�n�f���g-8�@x�e�t��o������t�e�V��?R�\ZVV�hC$��� ױVC�T�.�JO.����AV�fNB��{�ۦ�Z��ib��W��P@i���u��������`1���հr�=J;�ן��q�ܜ�����_���MЛ߈i�h���뫯m2M�ZA�?뀨
�ţ��^~��$P)h6AnjU����D�rd��#�&�vJ�ܱ�2��eJ/5k)����Ra���_�%�˶ƭ2�#S��nl��G����++8�QNC��|I���D���	�x�@ o�_�l;�m$u�ӭ���Z�e(@� $Q����T��.��5q�S'�h#���⭍�{���U�1HX�5�u�v�O����GN>���2�Gb�hV�Р����ȈU�>��4`�����@%���塉z<�"P��Xfx���
p�3L2ib)�d�y�G~���Y��ţ⨸{{T0ߩX	�!0-�T���F�S?6	&-{&�^�-O�{�iЇ��:��ג�衛{�QD�s^ m��?Y����aY�x��7ߓ	���aA�2G��e*b�I���v˚߭�gl�F�J?�7+s�;�J�ĝ^2K���Փ��
$Fq�k9�iӵ|oFS`��C6򲶫���X#d>;�܉5�ɩ��[.İ* ϒYԌt�˶W�o�cc$�C�6
���R�TN�K�U�B��^38�U��8��Tj��jU�(7t ��ʏlY��;�Z���uuƐr�P{�u茔/�\��d��$����}��tA�H�nq��=%Q����V(��݊��9�}��t����@��eΰ���N��K�#����T+7�a:b�4S�W�w�֣��B��?��g����q�H��L������.9PrG�Fi���nP�f�p
��.�J�r_�Zʯ۶A�<�N ��F�m�����D>4�?�F.���0nGRd(�)y�[�WP�����w�α�.0(we�7[Ѓ��8���p΄5���>3I���	�y�@�?>��PO�����[,̽
|���y�4�wg�%�����`qe �g%��z��Z�9�5��}�8���(��t��g6�f�b����]<^g�[���&G-8�h�g�m�F�].V8�S�����ЇC������-�F�Wi(��
���x�2���Ő�-ǯ�{�0;m�:��Ni2���Rm���N��rUI$������(����3����nz��$h�/�tf� ��}�~�BL�$�8�U��ù��܋�4�d���L䘜��8��7�<R�pb���%iɬ� ofT�ȴ
�H�1���ik/0D��
ͮ��;��o��N�B��=k�wZ�[������i{��+?#%yz��>&у�+�Ʌ���5EBIP\_�EUV E�_��z� ͩ��4��8��Ɲ��\b1�%�lPh�؛ī���,�A s��杖��&�Q�?;�:J��ڠEG�L�,��"��֕)i����y���_�|�1�j+ �&�I
��
wr,����&O��r#�R������v����C0|ʻz�]��x7�����:i�ƺ��(�W�X�KŘ�v����h�S���ڏ�W�rʡ���	VJJ���=������)`2̮��t����#!���'���W3p�@��렫W]������� T5���b؇�F�[;��qC;Y��4ߪ@%�����C� 4b�Ʌ��D�;�t 7.>�B���Gϼa�Z2�@X[��Z�6��������?��`w`nBԐ'y-xg���Q��҄��-h�Sf����L�%�U��Bv���`���.Î�_��7[�F���r/T��'y���3=�`�͋OY ����V��d�#�-�Ƴ���
X:ѯb�����qʝ{�o"9:�4Da�|��>|^!�
��:�	�x�f���5y��#��ot��8��&��S��p��p�cX� ��⯟-|i;*��?�u��}q��޳������L@���D.���ݪ%Fj���:It��-�]c�;�$�K�}Y*�Q�I	������7> �I�V����
j{��'.#���ݝ�O}�^���s�o	#j�]��sHFY��f�*���\��[і8���[�g=���fۼ1�?/�vؓ�PhR2���N>g�!��*Ѳ�7�??H��lw�8�Y&&�A��,1�
5�mՍ̀-�2ΈQe=���f^y�q�d>ɟ��oh��g>� q*�N��SB	yN�{h ��O�(��4��,E�#��޳�~��97�C���V��[��lJ#�#������*ƗX�D"�����ʟ1+,zHTSj��r!�"
`�R�� ���L��?�Ų�5��O��8��f����3J��N�so���~��5�d`{!((�6�q?�yV|��dx��{ԄF;�d����:Z�q$#�0�{�۷~ H0���V﹐���<6��2?�CIo�i%�m/�cZ���bz�6�@0�����q��4"P����HzB�q��;������������+�J�!m|*.�+hW<��D����OWD��qs:�ϮP�&�A98@����
6���p�N*R�>6�p�2��:����-x��I���{��Zo��0�׶=aŏ ���
�!\UK��J��"x1��@W���-�����֕���)��5d��E\�$�VI>���{�}�»y��X�5���>�O�L�o�E�&�%i��3m���QK�@��.�0��VX�OSgARH�5�����&Q��G���6�*t�Lu�jK��㎣M�Q*�E����#m���c�p: ����6a٦�����j:/�{��M�|�R�&���8����N.�'�{]7��q*% q��H�J�g3z���U������=���W%2�$7)z!��O�(���$W��m����ZgƠ�H��5`g��r�|�t�\���k]
��#0��N͌e%�)�y:��6��?�T2�M�͔W��{�>4
��E�}~�"A�y:3�ȓ��ǻ���}M����y�w�M��gU����Zd_{��ϖg��8� W�I�mth�\�I��}�M�a)���q��	����_M56r��W�җV�*	q�l�U�라x
�%<�=���c��s�-�+�u:�ƩM�ݦ����>	0�^8<EE��r=z'���5���1��]�/�����&IO�������/ک�L��<F���Kc�[J�`lh�j�U���/�XD��N��oo�.�
7�D�bRI�����Rl@)�Ӛ�Y�kt��b�aò���6�EY���F�ԧĜ2XL��v�7ž��RM-!���1��{Qm����=�PT?R�c�w��jƓaujމv�X�b��Ho�JA�[��m(u(7�l��X��9�+�
a��-�O�t�"�WC��XibE#�7�w�S)���Ե���M��M�H�������$�z�� �_8h�:DFAP�&�{�9��Ҹ�WCɚ|��e�يF��ݜ�H�����B8��&���̋�4�e���y������ɍ�<���}P.|�e�3~5���5ҹwK�R\X�2�dk���geUP;�,��.)(�y��_����IG���.Ğ�vr�d1B�Kr�t�8C[�!�TC��jM�=�'|��5(]��̚��&������rƦu3��9bo����Ʈ@Rj��I�a�J6���' �P�s����*����(����+�zH�lԠ�����K
��K�L�$@)a8F�̚��^�.U_�O��	e�@D0�a�#i�o�7O�X�N߹�P�5^��P���>H����X����h9S�6�ӗ�Àm|��SΆ�I�
#���N�]����}�曁o�Ѡ�uDJ/����ٶҞ��F21�l��iֆ��	L"E�$#�ϊ2�<��Bl��.-	�(��6�!�XD@�gK��bϱ��u7.��P�f�6��I������y4�b ggB�e|�:g�qq��Թ3���%��}K�<�$I~�h@���TC�o��On
j���1$�%8��@vErӎe�WD;�ל�@�n~^gL��O�ԮL#��M��N4�Me��'��|u#���0?����� ��)�f�,��沐VWX���qX�r""�i�q�|ǌY��N�:T�,t�h��/_a�͹�o��7�O���N�S�B��M͠�z �ٝ&�,tC��o�M�Y��XlxVHYEB    fa00    1630(y��F��G�.���1�p֓N��^�S�XɎW{��p9��rj��-vZ�Z_T}αn�Y�H���w��X&FW�o@E��2���8S����5�\�����;!9y����2\�uc(_�w�$��:i���~n��ݥ�8(�<�To������T���o��xݶ�G����zQ���ވ�?]����l9�c��Dc�����a�,~uL�y$(Y[h���m�[��b���"V�|�PM�Ѹ,�M�g1�%�_-P;裇�[�7��.&�՛L����Axq�K����y'N!�Y��vh����&�w�/Ƨ���r�RԠ�d<�A
�%7ol{@��wU��[���U�e���1.�IM͂���.jQ�!z|I9A&g�~�s������	�:Iz)�����B��u������]�믛�xV�7�{V�}M����g�(�^af敏	��|�j4h�CN0	����U� ѳyU7�*�0}�#6�NS�?���7t����G������,așn�̬㒺E���uWqG`CKT҉I����e�a�H�	0x1|O��`�".Z���۷,���:��B�ҔzM��<y�ߣ
�c�=
��j%M��5G��K��QV���ɷ��y�������r0��ya��\��A���y�ˮ�a���{�5�>7e4��-���KQhv �q��/�8�)��w�'ŗ0R��S�.�,rc�o�A���p��EN�� QX���	u�l
�P�a��:K���2zJK�K�!x,; ��l.�=���\�l���n2@Af!g�S��ُȜ�]�F��@���q��G�ь������-ɴ��R� p%B�N��;�Y ��;b�+W�M	�L�����3mM���v73�QP� �Fʠ*���b/��\�#c�"��.-�M*���2:{˔e�'u��e�Z�u�7`	9�Z�,l�86Ya�&|�%1�p��.��6+���l\HP#1�_v��	>0��z�1<��l�h�l���V��x���X���ˢ�s�ƥ�}�Ө��_��t����z#<v���8�Tp��pm��d��ϭ{�%��mXfĜ��
 ���+u0K���k��<�\*�o��4p��1�]�	�>�N-b%zC�G;(��Ix\��k������x5���9�pPcJ��@>l���߉@	��x��,i�~�͞o��Q�R��4���<��J�/U��N?*���R��#��f���Q�1m�4�Rw��=ۀ��,���dz j#�R��f�dΜ��w�$W`����uԠc:-��e?ⵊ����5I�U�t��+��_*�J� �y�'m���bHr [���\'
o��/A��{R�a�����p>�� �b&,w�`�T�Q�?6N���X�q���Y}L�ސ>I>z'�׉��>O]���XA��Vc�2��B�c�2њ���̀�_��
)�4�F��hM�$���،}�j-�<�ʷ�o��r�{I|'�sw�ƞ����w�N���2D*������''�|چT%�:�QY�������f�
í���#י@��-Fd��+�W�4!�N؃S�'�k�Ɲ:d�<�d����"3�{�n3K�^�ڵ�̝�{ �Tp��b9�Q�q-���w|5�U)�w��,�����#~ʞ�&r�}9&���c�Da��v� ��jߙ�C~ ;[YO�SZ��-�9�4oA)tm�j-�60����'�X���=� BI�+o��q�dl�aq��B��{����Ƒ��E�<�t�,�#��y.�F���wMe���-[r�!����e��R��:��*��K��fBƦ1�z�@2�Lh�r��M.����.�8蜑��P��jY�x�Z{b�9m���[�{OH�����a�30y�u���h+>w��`R��['.X�{���HmA+�	��aW����1�(']���yfq�h.#������4Z��:!����,�|��j�E�#��z�<���xO>�C�IS9u�������@dL��d�+�o��.���R��⮾o�]�~&��`n��Nk\-��Y�x_ؠ,������r���X���
�g�FRN/`�	�tIJ��$I�c��*��M��FG�P��!�3��@��`������Z�����%T_��ɉ�.��� i���wH����..w\8�ǔ)����p��$�]�;jղh�LZ�%�.��Z�o7��|�W�J�"0/#�W� l�������y?F�\�8|F�%�x3�y��=�?�q}��������|�v+J�1a�@*%�1["���
j���uH�X����!�1�F��Gx�8Rx/b��ye����2��H��<6%�m0ݬA@U7�hE�oa�{U�.�M��FE����'h�oo�Y��l����M�S�hdi���e9.�,6���-��bZ�<�DC�r�$�/�
[M�rET�IPi��b�+���^8�n������#�ù7���ҥʨ_���{�T�>̒^�r���o���o�f�N|�Z���>�j�_f����6nb���|$�����Lڌ{����u�9���hXq�!6Q��,�9���d�]������Vn�G�d��Gӓ��V�J`7�� ��5�C�K@]w��Y�F���eV��-�`��c��D����U�O<��#_���*�,E������'�Q�v-8-ϛ�K�$XeԒn�%������핽�7�ƈ�N\��I���m��ݯiRˣ��Vlv�h�sZ%�(=5���"Z�Ĭ���������Bvڣ�8��B�I��a���S�[�d���`B��%�"�dh%j3$��k��ǍA�bY#z�a����dh]>�3-��3�<v��a��-j�aƬrT�dj��&x��j�t�%�r��O��$uJC�y��a?7��t�抚"qٞSB6[��e�b�DY��ҕ�e��2���v�Z��[�X�bN�d=r�Ml����m���:���(���_J�G| �]r1��#UG_�.�r��e�?��Ɯ�&xѬ�� +y����r��]M�P4mvc�E��J�&Hӣ^�F��(����'������^�Y]yM"-6��߭��ZQM�0z��r�Jh� g���ǘ��1�`~�P�!�j+1���2�y?�8����ݓ�� &�Z���.\w_
B�(|�z�g�hR\:��I�a.�k�(6������������'4cߞT�5<���7�?�Ј��x%�A��K��3J�CN�2�Œ^�1�o��/Q�� ����(�Fy�g�7k�fʑ�JG�:���GU ���%\�quy�Hm���#����j�M<�����=��m�:$�J��M$����=xS!7_�7�őQ�~l�`]����/�ܪ���j�<��8�&`��&�0ܚ��n��y��֟D5\�KtI'GT&�_���JQKA!~�u�t����O�tK;���j�E����4v�w
V�!���9tv���F�swoԜ��K�P�������tdodc͈Ġ](vi��0I>�a���-�����}�׳(~Ӥ!������F��m$�)��c����Ga��G���cp��㚯�>�D[��0;�xG�1��mn��eb؎�zT \�:�����c��@��7�~Z�}�b�P��zJ� �]��`�P���va�����Z����7ƭ������Y	Q?��v�s�3�>F�b�C�=Po�����g��xɢ�Ij��<�5�IK�(R�Ij��?�Ǐ����W4	�H�;�7s�����ֳ�j�I�X�4�E3�A��;�5E��KK���]����J~���+���6����i��h�4��>�Hl��/W,��G����21�9b�z���7�BWcݫat��[ޤth�Bt�,<*#�Vx=v�KݻQɂ�`�#"` O�4��i�SQfT^���0��/�L{xuRe��x��&��
VP5,�NRƯ����MU�]1�ψk �Y��.���y�>�gb	��^��>�i�I(1�p�2#�O�/Y�'[���,+�h�}j���5os�4�$�.}�;�c|��o��n��]�P�[_�2���R�,�d�x���{��=�IpK��څ�Q�B�ym��a>�)K�K_�ߝ��p��%��h��@�5�S�cg�t�8��^�W�B�։�����׊h�Dt6�8^���u�������=_4~�,r�p�V+" �9ɭld���rq)L�m�>��3!;�׳@ ��4��cM���T�L:X��*wU��>����) ��/'�8���Nwg�u�7�+ON�XԢB)�"�ԉ|y1Y�OƑ鯑-`mAt��7Ƈ]aܵ�	3�a2��D��r��˱vm�ol�RI�EF=�Q+�5<H=T�Y�G����)+drl���_eC�26�YU��G�H�U�,�>�����e����߯��:�ѝ�b����d��^yk!��G�:�:���a�҉�:��c�3���C�r�՚{��ʋ���S��h�Z���������w��`^���[:V�w�h�9G����KR� ���Ǽ� �>i(B�<^!�lq'���S���a��Æc�=>F�<x;/.���y��Wl�G��J��O�	{�GQ����G}8������(�h ]{�~o1�ix��\ʥXt��!�V��=BV~ܫ��脖��0��l��,��dKp�uGca]>Z(z�,�L�bp����ɋhW��Q��0���r��������j�|�LExְ"M�߂�ܣ!�ת:q2��z�k�bh�P]�}���J�H��n��^^8��W>+����В?<�R����A2��6󝓫��4���	�Q{�d��������e���21u�H�!-�߮j����3����c�ޘ5���G�/�e*��U#�D=���9h�]�I]�\��<Y;(S�AR�n�N6���	z�}*o�-��m,/ȓW����"4�!H�?ń��<H	��Dw��?�q�fX$�ƺ�}g�~t�tꂩ������+~d%����BA0S�vGAw�G'��M��/��@-���`͍����ǹ�ix�4Uۦ�:R������
8?�-s*&stΟa�	��ۿU�?����h�.�/��[+��L���vJ(�X�W
����a½�o��n	�ƞ0&���vJ���e8	G�/��Y/��b
�b���]��g
Fl�(Y�"�Ѣ<��q��al�q��_�9���a�ԁE�����0<?��=�ߑ�aa����m9�jx�a �c���Q�J��\�[̀��E����<ǒ��2S�����Jգ���hu���{��	\Qw]�O >� �X���񱤫7��9����q�`>J:��pG�Jgj�j��(1���o�H?=���O�d��2͙�qY��,�1ux�w�q5��I�"9w��\?�8��`���W{������ă�_��E�_���fc��']�?^>���D`��'���@C����i��r�LD�,�Ŕ�}s>��p���VѦ>�{�q̓K[tC}��[ L{�z�"]t�z�{�oZ ���H�me�XlxVHYEB    5a90     850w�۪d�Ef�*��ض��'!�H%z�]�i�uR��o����mwK{��E��?��S�'L�J]R|��j�\cbF��>��/�S%lձ��;�>,���9<8�c��^�����a��tx(0ܨ@Ȍ�^y�JVP:j;���T�mLrl*�����~��\�	�D�ۄ��z74I�-̍7Ql��}�,�:�+~���d"�-��B	��|�|����N�7��qȼ���ֱ:�<:�G:�{�Ԫ���/�/�Z�z�ޞܖ:AH��i�����?�PHz�����̜ *��ώ��@�#�7�������ͧ{�Q�v�Y��TN��l����6���(�@lIu����������;ř�BL\1��EbR&_{L�S.�y\o��%�(�Th�XP6�-����;���JqSi�#��>���&�5 pߘ܁ɴ;�¯�����ڐ"�7���EZ�ֆDi7��9����$GRR�_I&�O�,���$�#�
YIm����4�dD
��c<�-�%��D�A� ��x�����̃J�=Ӟ�Z&8�9�B#Bk,�Tp�m��R��d�pe�G�P�V�x�:�p��띚���<��`U1q0l�BY�D~Y�>I��R���Y���0.5!�|�z!Bs���EAF�Ž9�-�F�9��$e�]�7�x��v!��y[���mR0�:��>f��~��O��_e��
���Ӑ�@j�Zk��:��+��e��{=]He��пx?m'��� �d�p���to�0��,��:k��v�(�@>�b�ۢ
Gd�G������Q�Ga�Dw����ҨBӴHq��Oǘ���TXOl�-�T\�I��n�s�Y9\7�� _�	�tE �<h\ڧ�����F��u?#�fa��*�a{�B���I����͒f)���댲k\&0Sւ�̶����-D�Z�Rꃿ��&u\�e2�<\s7ΜM���/�ژa�*������u�;J�謫��DNN���ڂT
6�l]��e���6�����B6]#c�MD鞩1E������*ԗ�q�oM��d"����"#��aB`\�����s9���_���6vʞ��7�-�Fv��LK gk�_�7�SE�b[ʸ�fO��	\|�|SYL�$g��j�@�S�ʉȺ�~ZB��/�\���'�h󒧻�ꔙ�w_�i9��w�$^�u�X����+A�����ē�����a�d�����C$b;Zf�M-��PM���yV�Wkg�kG�ۦ�.^ۓ�G�wrE}�_�)�1���4)dޟ�K��FO�Jk!,�F�J�&B��P+�����M&2���dZ=�#4R���>��Y�7<���ى_��Ǡ�<�X̹96�&�h������0��Y@��]^�e+�Y�?���pmz�g���i�C�@��t��y�����kt��c\ռ�w�>����u2#�_���ˀ��"
+Qv/�HD�崉��M��$5�ȭ�0Q��`��7�bU��$;�aCK�i�Q	[�"p�>|���w,�C��rp�G���GV;v��[��/�0���ƀ���_�i�2y� O��[�)��	z�����R�> ���*�q蕦b�l�Z�;/m�/B��@�������o~m/�xĲ#�9[ĸ�ѲXM�P-�?�����̬oڄ������癆vC�/�6�s��2'��b�c|�2�&o���S%���S��EC?n4��܍�uk��"���u��'����$��F|jpa�fW>~È�.H��-R�6��V���>��g�|�0u�i)r��=�,e���J���᪬�De�������"�C��	@*Z�i�/���&�jk��@:�u�8a��؛�������Ze.pn�����G\��V䫑�j��~B%$S�.b"D�d�_1I�!�#U!�j_Ȫ��ǡ��W�Rg�Gנ"�ПS2n�m�P��@���;���� }�1�r��a�g8���Yx��Z�`nM�$a 4�Ϲ�R�z)2�s?�ï�*�9�q��-�)8��8s(����4���p��s>FIF6���eN|���]�Q���91���:R�nbDhg�%��