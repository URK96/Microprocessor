XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����{�=i��O��j��V��~����耡�_�\ў��P�'z|��CE�]@��$H��ؽժ��Ev,Y1�`S����l�ɛ��qcg�$o�*�>�lwR�,?䲤�5,U`����js���"�tӦ�8`h��M�b@�c���@?f��Px�*Q�y��#����-H�?��F4=��I�t���!.m��Ag�!������3Vu�/�om|�hqnZ1),���/�D��4��<�BK�E��L�C��ȷq���^
����}B>j�50�m���#�}d��k�B�@��e�J3��#�����W�?H|h�O�;7u�^Y${
<�Qu<��np	Ovd��9����,�m|��v�c}Is�������^���������ƚOI����*0`�ЪΫ�46�*v�Mq.+k�����%�����/��.m�e�!c��i+ERD�þ�ɱ�2�]���OqfTV���ӫ�Q��:5ы��B'x��h}CE��d������3��J���+��$t�ڞ��`�H�a�\��5��>m	�ӂZk�YI��@ Za�UP�]p�S�D%����ĥ8��}�^lF�uZ �!5k�A���8���D����Ҕ�2x����Rs�imTko���~��9>%��R��_�za�'z>ὑw�Hθ)+�t�h�L\h��1�u� �
�,�A��������MI�[�B�;V,�CL�Q��Zq���s�����<�9�*��hB<��{zSXlxVHYEB    1044     4a0���AʺwQ|�'q��_�-���b������С�(��!�D�QLnk����Ƞ����[I��2ۈ���H���$mZk� "w3z-V��>P9�vP�aW�X�nT������s�],w��ҳ��nb�ZAt�����2�#6��8
~�t��!֕��sJ����Z��J����)q>ӧ"������"�Spqɡ?�s�;n��S��9jC����قݭ�@���|��L���m�H�����Bv�ӊr����m�y.2v�'�X��e �d�l�HW��u[%�; �=|���-�)�&^;/2i�����*�&�
�H)�P�P��T��즒%��T򁀥-R���p�Z� �X���n��]_eK�(J��Y
wϘ�FL�b���ue� B�^d����uĈ�Vn-fB&`A�.���/$ȱl��1G�O/��i,> ��Ҙ��jw��)ح��إ��R�w�A`4&�Q�;bB�� l���iI�O(oK���@���*hv�g�"9 ���F�vCJZo�ّ�d�ϳ0Ʈ�!�L����JxZb�p6(���\őU`s��h%�������3���8:��]��gU�& ��H470�UU�G,/E�6xA�!�~��z4�T�$�sz���0!Ӆ�L:2����k�?�!+������Y��(Xd
�3����Z���Q	�a���%`t�=�������E�r��,�r�E(s�@��1��<e���A{?3Oe��u�2#�odĉ3���X��R#�xku�y߂>{-����Z���!�<O8�^� �t�c.'E�ׄ�	�'���ɹB�������ǔ�{p�6x\i_Q��P�ݕ������ɏ��~�ҋ�٣%����鵀82
}uD�7D`�<�+��;W�sa�:3���"��2 �]���3�-�BP���t��S��!��N��`E�O�@�E��/(�E���=��!�ʢ���n_�y���u�Z4_����]�]�<�
m����I�1�v����&�����)��i�ͳ���GA�1 �B���'��1��\�*�s�g��LDl:R�>�����ضDK8F��6a����nh�~7|�}w�[��|���-���!���I��j�+�Xh#�dY�& G=
�(;�U�z�