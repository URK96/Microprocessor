XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9�m.O�:��C=�����'���.��]<u�=��䐹:��_����t�o����Z�(����^F�I���i<'.}X�f��F��^��m���:�8\��,v�%�����"�� ��r�>d��$��e��n�=d��p^�D}$9�s5RS\�F�$��bP�!F�p�[�//n��m�C�q�r�4��'�{%����!Z�	����〠u[�_@R���nc� �M[ЉoXE:c# t�eK��o(�_����;"nb���%G�a��%�V�nLn��ުjqQ�]�@��6�,O�aԓ[q���3����6��z8J���8GT1�ZztP���E�\�җ�b�?���^sB}F��۫t{x��JTV��^a��3��\v#^qH�xq��3_"�`5�q+"�ښ�X�j�jc�E�k����N+*��;b�:��%���gb�0A�Z���f��,A��T�A����9���l�1�
�6���^n���JD#u��F����ˮc�a���,x�1c`$�q��i�`V�]YqX=�_m<0���փ�oP��`.:h�mx��M��;���kf���3����9�#��j���FӇ]N�IN*��g�DZY}O�?��_�ִ؛vc�ה��f�.j��&�uhU�p{HIO����׺Q�~"4O��ڦb�p�x5��oP������ �~�EF���R�ԧ�LX^w	Ӱ��d�&K��V�L�^'��cE��?�ٚ��*'�XlxVHYEB    1cf5     790��S�G��.��3�}e�+|N
�7�/i����cA����;8t�"L�� �/���w����0�[]�#7ZO�߃pzi�������������h�iM&��`�$��|�u�k"��1.��G.J��F|��݇S����cx�6��:���B�$S���y�Q�jn�Fu�9-����B�s���^�����c�5z��5gwזqu�S�l�T�a:��Z~��m�j;�#��L��D=��&��A���=X��a=�-P��QB갔����=�LtXr�.g�`����!-3�f�zG�~ȡv�>(̨b�+�
654��Y�4-g"w?�d�]UY(� ��P ���)̕;�w6��-,��9
d\bV���=�<���; i��پ��fG���|�U@0kk3ۼ�yR>�f;�iԌ���-�y�r�?UC�j���uh���LZ��6�ݭ[	#Zo���h���q('����&�T^��nGĸޜ���Wx�pYH���t׍��J��K[CFV3Gˈ�n��EzQ@��:�lTnq��4��ߍ�W�ѡpN�@��A���C�K5U8 �S!����h��:����������R��K���5D�?��#T�ۆȹE�����R_Fk��u�AH���6?k���r�3,$`'����|�x��q�@��xΒ_@4s��#A�=!�s�� �`Z�I�q�''"�L2��@��dǉ�R�^�,ܔ�[>߻�I�!�*��N��X�nA�g�J#�ap���/��(u����T��=���.�`���d��V����G �w�I)��$G��)b��Bc��V�?�F�xƮ�/�Lz$Qr����[@U����8������G;��.|�)�
�8�I�Ճ���/�B�A�� ��:�0��yʔ�ؠL���"l��N'Y՚Ǩ�,ȹ{�I3#1�o�?_����
�e�+:d�����Ԁ���8������eG��f�h��Iq���0�-��l�i8eX���!ٓ�S�LC�FQ6�R	��S3�W����ٙ�N�C��`��U�^�,#�g.+��_��5�8�s�Xtc�1=�Nh�Bi�%�ck}Dt������7SC|s&n�@wr5{¤t�sG����\����O��*�U]X�e�E`�(�8��顇8�.��y���y�U��I^�|�z�tEV2��T.s��Sj�N0�m
�z&ks@� dl��x9tJ�O�������a�.կ%��9 =��X��zI�Y������
JMZ�	
�r_�����J��ÏY"��N.�Y��M���!�ۈݗ��dy�"1���i��ȢMIأR�n�փ����Y<Z��]m����_��I� ���$���NH�1�֋)1v9�ge��?�矉v�;)���.�
��.�%���|�ʻ��p� ڀ�z�sF﮳t@�ĺ(®ƃW����d��Gєߌ���k������,���'�s��T��[���D>�]��l��m P�� �>�;��QC-N��,��j�����f$�-1�¢3�����xJ@g�������bȡ4�d;6w��"�p�Y��WBj��}F�U�߮S��=A�aW���+Fp̞�)�+	����w�504�/��>;�,���]3Z*���m޻Z	��xvM��O����@hύ	=���[&x����V]A�Q��h�����A�jؓSO;vM�>rR�"5������,��d��Θ����)�Ć�t.�`p1Wuy?�}/���@E�uN���V.L$NYQ9���ƨ}'Pxs�h_�g)v��� i�r*%R�J*J��-�VG�@��]́�
k��s��R1�MT|\���
]U��SdZ�����_��@Yz@����\�yl~��Xq�:L��+�N/�WM�o (.k�_