XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��M�V��>�"M����#6��T�QتUϦf�T�l[�S�V��X�`��N=�P���|�K���^L��&"�N<�G/�X�>E�jZgA> (�ȥ�bY���lA�����8�+E�>���霏�(�k�񜐊��a�_��B�
n����o���b��f
�� �M���R1�c���^m@L��~ID�X�MD(�BF�1`�m}���s='����H NX�~	g�#� �j\r��킵���LE�pR�-� 4G�i�P� ��҉4�5�:局.��5�p,Q?�Y}��*����W�%�j_X�|X6�.�Q��oOJ�-�0�Dd�LWi:ӱ�&#�0��IbU"�1n��<hYu3c �<8N�e	[��,`��j�u� T�R�٥���#g_M&ĩ���M�4��aC�d*(4��}��um���F-�,/�V((�?��D�ƽ\-��;Ox��FF�FBL+�Iė�����A��՗|��`����"��1t|�6�J��d��6��"�%/�l
��S����a���q�1E�g�/�!��Vd�m�]X���B���%Y?�f$U�W���r�Q�u�U ��b�a��m���K�_��ז��)��:`b������j
M����L�PFV�4����Ѹ1�}�l<�NJ"F��=�h�i���Ǔ��W3X��C�� ��I�T?��ތ����xs�s��«��a,�m%��-kc#���БНҕ�(�����'0@��XlxVHYEB    78d3     da0��ɻ�p�w|`>`�̯3U�d�9}N@�\lW�L.=�lwhH��U�`|
��D����"�]I]���%+W��i��ܪC��A�mW斬�"ZTF��D>�oXu���DEѶT�*����/��|1�1�a�ŴYdt�:Gr
�)�W/xf����#6��]B����(S�3A��`��V��U�����(�����FS5�k�XEN�TB�%���#c6r����T�';�6�7�pB����}��F�Jt��83 s橴Ak�������J`,`$��zF���P�� �?BG-�8�@:��g~w�;������d?�J�8\0ۃ,WJ�տ�Y�z��.�j����6�:��!!�J�pl�Ѽ5j:c,���v}���>�n_�9{��jj�j��m��5M3x%ܡ�&�F$c:bz^C��s�}�z�����W�>���ҍR�����ΥZ �4�OrI��7�Eb�,�_T1vZ� ܂�tl��!�UH�]�A�:�6\�fэ$>1U�o��<ō�l�N��n�2��DІ�ѻ&h�G��	&��!��3�p��P��D�b�l�_�Ƅ�q��:^�\�%�c�kG�v+9�wX�f�R�q7Fj0�\V:�<�2i�` �S�贃̵�xK��|�"��3�����z����%t���2VZ��g�\P��$���m9�N��lv�������C�S@�?X��q����t�����{ �R|�^��!9.0�BJ�C�[�ڗ.߇�hճ��Gv������z�r�tX������H��'�+E�L�}��J^�CI�Li��ؼ򤜭6%a�M/`�rU��)����q�������B�o�Tj���8P �p��C�0+��6� $� �aO.�ރba��hT��!�/�U+ D�Z���PH͛ks�����a��@����on�a�A۩��p���Q���˵� �����k�����U�>%���!�X�yP��s��0�^ho�5XCfǬ��L	g�q-2=��$���vԙ�yNÑ�'_�-ʮ��t���_�gz����]OhN�@��(5�I+����І�����~I����r9��O�0���|�7P1���5E��}'�^5�7<ND(;�+��}k�R��F�GnF*VԀ7'eP�zIa��$�xO��(�Q9�FcS���"0��!����Lƥ�ix���s��I��K��['�|����C��}>`��5N1 Mvcr�����%^����3����=���w
�F˶uv�ba����b��*S��j�����o����s����HM���B��@_�c������GQ.Ľ���~�����e�>VS�ok��E���P��ǥI��L�`�H���b� ,�R*V��X&2/�ǩE����F������'�6~q�Q�4��H�
Գ	d�L��vV��O��P�Ҏ�8RclR�#�&)G�˳$db3>\�'�G�sܰ��jךf�2�Wh��B�R�O2�Y�&Yw�t�P������d�r^�T8���#�TvTh�=J����+t�׉c��3n��XRmz�Q�%�1��6K#��x�������	<aΦ*Iʸo#��fìIqT��MoO�W��w�,,�e� ƴ��<�<���˅��x��Ε��R����d���6���S�u�z���/��ο�
(�
��:�����(0$� ��E@ׄ��eՖ���<��|��"���}v��4!85$�Y�]u�d�9�pãe���X"�������Q�	�a�y��	�{��At�� �6�}B�&����dG�h�%�	R*ND�{�j�z~E�S7�8�4�c2:B�Er��,)[��x��KH�]A�FE�20^+9���:X.L�>�3]O7+�#���ޞƈ��fRφ�I���z�NÚ��ڥ���
����8X�T:d���rְ��=��e�3�gMB�'��uN���H��+0�Eʔ�	;�����kER��N�75~�	*0�WLH��Lb�G}cH��yP
���"5�皥��m��>J��p�$F�X�*�V֏��^۲�25 3^���5b�0h�9|�9|�8����@��0��!,���`���g~�i��U�~�!w�)�$v��Z�b;nU�����e�{���MT�q�r�/j-t���b��<j�J\���������[�q.�pd���~����kJ`+���n��r5��?�^,����׾���zܥ��C�i{�ӣL�ؙ��y�����k2�e-��V�#	I&P
��P���]!<Sh��7�e����@�x~B��Iu�rZtt�<�#���0�;x2n��Ŏ�U��4Z�I*{�qС��n"O�;?�0��`l�ŐK��l�'��hR�I�:�h�t����/C�k�goG6���u�� ���s����v�<�ě ��R�e-Ϛ�u�t/wv�3��D�:����,I<��ݥ�ϲ�B?�웗��q  �P��N�*��؇x�9J����2y���/��Hؿ�K�d���Ė��:>_9�d��X^��%K=�q#��!mj�oNR���q$�],d`��+�%����8��U�a�qIoQ����|��;L~�jl�Z�����/B�6/���!���;.�f�~O�t�c�pE��o�C��1�<��uRh\bYr��EL��� M��ifyF oa�c(���B�ɪG��N������uR*mz���Ioxdڴ����Bky��/��T��6��}�,��ng�<ccG�Nx��î݉CMؚ��r1�<����QYt�Ζ���`�����b��,-�����������OKC�磖q;s��	2X��L�����c�'��Հ��<w�ن~3	�e�>:ޏ�_�5��iA�'�⊞��iٸ�I���9MX���L{���x;�ǵj�(��ġ�S�����Q*�⑾G�Qʆij���M�]{�ec`֎：��)�%'���-�T�5 1���ú<֥a�V�_�39�������u��_KwMz��
f��ޛ�Q�M�q���Zx��������|���!��#�v�>R��ঀ�(��Jd�.*ƽ��, ]h{��
�{)fI�Lϙ����[��b�ϸ����؈�]L⣙'��N�-����_����c��-E"�w�[Ol�\���w�*	�s�~��s�k�X��{3�۲��ߔ�b�?IY��w�ee8���w7����f��*�zm�].�;[�I1ENA��ψ��X�}���,$��T���Z"��"��w�o�f���%c����if'��Z��P`T�L�cd�8�Q������3nd�mY��w����ۺ�p;3���"B�y�i�ϣ��g���[��t�Bȫ���Z��[�=9�O�oѮVt|fAG�}�K�G�w8Qƪ�D��ic9�!��bb����u��,�Ҷ{�p��R( Z