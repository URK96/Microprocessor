XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����;��J�l��/��,]TfRmIy)Q �/����w<��A�$�ra2ʦ�y�F]�7$����uOgu�i|wa�ea���ȡ�*�\�**X];��]!�3v��	�ˉB3�𓮌����ڱ!��L��kl�aij�_���Կ�1s:�)��Q@��.��U�����Ѧ��L�"@K����i�	B��%�`�E�[niI��2)�\�x���I<�|q`�a\����)c.
�K�t|��ɮ%oC�A�♃I��B��̹h^&�w����"�_Q��6�4��ۈ��ϡ�z&Tܣ��^�t<�[�t����E�cОW���P��M�O�AbMpn�!6�n�~�Ws�~h�b��/��L��"�h���3K��(R���,�#a&.j�����#��LC��A^�9Ǜ��1scy:;v��Ѽ���)���a�t�6�t_�IpLt\���3��ܛ8�P��V��]�;CC��n�puH�+�����8����N����3K9j�(�"�2���W�٥p��<����Y�����/P�0\�F���#��j���)�au�Q4�`�3us��4a�uEWa!M�j��k2�2%�.Iq��@��I4L�ʩ!s�����'ő�u1���ځ6��Y�����k�845>���8f�GH���ﯖ@Q���m-%dq���J�]�������=d��M~j����F�����8�»�>�)\���6�������.���x��0�w��b�|����S�����A����e�{XlxVHYEB    3c92     900�MP�R5/q]u�S�2�ӱ�n0�#~�J{i�F��[��RQ}�bs��]�l�RE�o,Si�6�|�Q� |�B�f��'�*�j�2�ҳ;�}\��S��Mr֋�U��M �'�M:��R��xM��
�u{�E>��w��h3q)2�o<K/�
��m�%�6ǟx?���������9�HW�OѺ��g7����1̀W����~�<r����	����W"*�lO�b�{�T�ӭxvl� �H4�U/��i�ѐ+pY�3�U���d^��p��BتAD*�%�_�X������l ��hx��ſ��C�Ce���>�x$Iu�&�/H�c�8Ǔ�Kh�%Id�FBD���R����9H��bj�=.�ϲ��,jJ>��_�ߧ�G��o#x�-݂5�Y@J
R�����Mx�s�#(Q��l�YN����R}�������p�@�Hxt~&�-�����o�趃*7{�����@�
37'{-�a����W�߇A��'z׋|~���������k�p�N4����7���Ur�-���I���?Nk� �K#��j�s����=�3��)�wL'�Ή���߲o1zD�jR�`�T�[��
6�f,�ݏ��M�J�Ų$�#j���1�g~JX�<�Ǯ덽�v׳��Ĳ�. ���9X|��8�@�U��!�82U�ۀ�j��<���>����R�==���G�+Z�7]�h�-����Z�Z�Pwx��J�����������UX�I�au4���0�(Z�H�>��|�=�� �;`�%ѻ�(F�'!6/P?�<�E� W�4�2ȕ���]'td��ߧ& 'k�B/�%��܇4t�+��!��&��G��G�Y�g�h�*���Yb�y��5ą����nF�u��ĝ��{M����!YV'i"�G��z��`vj�]?:C3h���30�ч��t|��G³<�u���۞d��W������b]���Ʈ�F�}u$��<=�^�9e���5A�j��.FFv��&�?b�{�g�[Nߒ�o"}����
���(,�ĩ��Y:�ŧ�ň'�4qd���@�ķ� C���CXb\�ft��v���	�%W22��R�$�C!�=_!���rV3�#<�x�=j��
p�]�{Gʬh�b�ge:Q��w����d�=[��e0��Y�@o��G��6W>�����8����C
�����@&�,	�pT���DO{��E��O���^�Et��pDÉ=��W^f�� 
'h�#Ҁ�ܲP?r�-^�e`�6N�»��vZ�ϑ��c��#Om20��6ϲd���oT�tu�{��(r��O�2W7�� �s%`�H\�B��M�-U�=�_�i�~��߲b����:��X1M��Zt4g_�~E�:G9)������I%W���^�L��?E	��C�x�f�;��s�-�J���~+�=��+�QF�޺�ğ�!�}g��B��Ux�̧��2�~y05�"H�ӛ5��
\J0?M�'��3Ф
��oW�y��'�wUt���MYL?�5�o�����v�n�Cj�+x�C�P�?�>��Fp�
Ǒ����T���?K�������Q@|�ш<�N�@h Es/&�E�q�\�[�C�f�ڶ5�pRF����-�|x���A8MQ|Nc ���m�dxˁ���<\�|�xP\�����)sy�Ds�ApW���g7��ky�c�*s�H�����ž��?�6���J�����g�������*'��.��W�͑X8�G]D�r�B�!�av]������)�D����:�\�#��{VU�{���"�oN�lD;w�Iq��������v�a���NfW��Dbe�� 6��<f"��#�?���9�,Z�VT�M�x�xـ���:JQ:(�	�\����(��n�K �bMش�خ��I5������q�r���ؠ�f'>�2��[��V�	�
3���0���|>�(ϩ�<9E��ѯ������Y����25�J��G�5T�-�H�µ�
EOsM����..�a�ay�}�k��6��!C�<�q_l���1yE�K<B����j��a2->����΅�����#g���ݷ}.4���}�y��D�?+�lT$ '�������Dغ��r�H��T0p��+�?*K�[����h!����Au�r�S�e�Ԏ!��Q�]�&m�蚡�pƷF�x�CQ�����(XJ�d�P�߬��D�AJ���"O{�;8������~����NPl���b{3B����