XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/��^��6{|�$�[�"�FA�`8���W�X~�C��}�\�ʛ���!W�.�c��$䧝�ж��I� &*O"
'�I�S�;���Y�M����$I��@$��{ Z�R�R��`��eq���:U�h!����h>�&J="�inB12�#��K��l ��5r��핏B���K%܀��	k��r<�H'qx�H�KR��F��GF���[�v�톃r��N;��#O0q�E�bn���4-�j������	�Yu)k��6,�p�Ο��3<ܚe��w��W�
�x�����������GT*w�h��p�>r<WL[׊�#ct�}���ZI�f��ҕ��͉�s���zW)�a���d"{�&Hl�)z{���f�pk SA�)�qܶ&6��vL��\��z}Dt�ܮ����`����9_�O��������ρ^yEg��Q<ZI.���l�v޼��g��Xe�(E ��	�hF��axo'k�,����o;�[��3ꓧ]	<j:���}�(�D4�Y��z�Q:��2�,Ip,M�b�\��}�;S�m(��#�ۖ�Zpяv_��V��Hַ�
��1�"(�Ұf	��3���0,U��
F\�"0��U[�8t����u/���I6��	�#�%�:��<��Hp���P&,��}�c�C�9�����و���*C"Yب\�;�#��+�v[�2�=p��R�-G���� 9�3���7V�:K��l*O#=�<1�?�{���#y}��͡cke�);���XlxVHYEB    1046     4a0�� 葒�i-��2v���d�Oa�#�C$����ƅr�v/I�*QΏ�=o_$ϙ���j]�����z�oU�N�i�؞W�1� N��j?��Ƃ���*�~�E0��QQ�[��h8gݽj��w�<��˜�:��J�?�H"�}��YG]�O=���'QEM�+N���(���������
Ǭl�\Q�V���K�WP@Z�Y�!6���u���;�����ba�7�2�俐~g��&�8q�Cy3W��<�-n��LM��cȣ�_�O�oZ�=�s���K�F~��&?��ܢ~�Zը�D����11ϝ���d�eg ���d��� ��yѢW�k-���+���9Ͷ?Ju=�R�J�-�s�WN����k �>~e>)��	�E���ڶ�\X��~9� �85������'���oz�����&��,Ɯc5�`���vI�X}Sހ�Oz�mz��t���9�n����l3�G�Ed��$�!N�.��>�ΥG?M�q�|^R&�"��,�k����n:ҎP�Y�jdb�CY�O�f�b�Q�5���"���6beuj��x1'Dd>o��Z�)ݶ�2z507	죈G\��ˠ3�=�[8M�网��Y�X��G��-�C���VTs���l���G����,��@u���E��i����@R���x�	���Z�� r5:q]E����zI3�R�#@�Op����}����It����RH��O�iG_�<=�������{���wB�	�YjLi��zێ��Cp�W1z6}:�Ƀ�r`���9}H��L����L�Mb]����z[LS�j7�MQm	��^�a��]"ۯ�5��b��.f>����N��٤��ѹ�g�4����= Ë�{��s�T�/b�.�8���x�8/��Pc��S拸1����S@�!䓸�#k4��N��:I.�e��gz܆;����Szs� g�'e�𰢙�� �1Ytl��46a��pO��i����IU\a�rhs�ե����H�?l�{�Jx�9�Vt�3(�no����.�\5�����{�w6�wSǇw?�W�õ�PC9y��,
NsA�$9Nڃ���	 ������Wy�2b�����hk.�P�oҋh�~�l��t�t3So�2�,,)niM����