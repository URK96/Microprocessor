XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����J�C�����@]�#��]	%���_"��C�d�c�Y�w�`� ��N�c3<��Q0�U���qӾU�.�2�g�s-�F�Dp��6��f�(Y��/��UȪu b|�FՌ��[�22[�#��[�ʠ��>�K����^��`���Y!=���n|�	��o�޴�(N+?��8Xl3�F�	���۫3��HR�P��{v瘳w��uSB�6.�(��5*�	��gS=±Y��S�9LM�(/���x�F쇳h�5QU���z
�(*p�#)�>��_1��j}=��px���k��hjc��s�i;3� H��	��o�Ʋ錁�R��Qy�|_آ�I�.����RJ�\/sM<���䕙vR��"�`�?�k��	%��×��R��=S�+��͜%�`�����)�(@�{Y}X��)^��P,tj󞫰q����:�o���R��3p�"�K5��Si�;��X�ZŃH���������e-��5Qb��5�����Wh��'M���s����v�|j���%�i;� ;BZ����~����Kc�~�G(>�����BJз�|��[�!��]��F�)����Ժ�A/.:�EBj�=�.���9�4j�=}NO�)�P�����6�g�9ݐT���X�Uo��գ��}�>~w�U���6��M-�IU��UՋ`"�xL
��&YD��jtţ�E�Yv��F����ԈH4����N�F.NDħ0~H�P���55���TP2�b��F�7d�W������XlxVHYEB    458d     8b0����rֺd��+_��+����ᇢ�HϬ���0�g�[.5W<�T�N�RY�%�zү��B� GK�";�+q��E5!ø~W�p=|.[l#d�F�(j�l�3��������	�͉��&��V�[G�w�2�Oa�rc��Z�x�X;�:�EC�(>�:wJ��#Z�%����	@���� g��fvT�V�`n��Đ��Ux���d��7%��d�/�Tb�4g��L� ��; #-��x�Hv�=6���Z,h �O�,O�K��,l�#��j��T��S�u�Y���ܶS�Bjμ��Ҝ�Ni�G}��m"�l!/�J��Բ�*�&W�5=Wێ��y������7~SO�X`?v�/f'^��\�b����8��̾ǝʅ jy��,[k��C�Ot�K�=�9�+�8��y�.*?CYGT(v6�Ȟ��T�m`D����
��Ϝ�y�i����}4>gϻ(�� ����YI��4�����t���j,�J{�=�k=�,�4O@S��0���5����	i ?R�A�|
����S���m{j�\�G<�m ^��P[��a�����'��4�5͑[B�Y��������5J��2^ؠ���-�ȯ�i���l���ȋ�o�6@ڜ�����tR�΄𭡢F�gp��1.�&��9�oi�T�>+��{̬� �'Ӏ����Y��9/޾�f4�������G�P}?6Qny1�át$%����}�|����9^^Xu2��@E���j�=x���ݾ���0.(�C��Iy�3�PXI�7Tv�x���;d��ib������h��&s����J�Xl5��\��ܕ+�im+�9�}d[~?�˞
��6��sےʉ�e.����_��Y7y(N߱M��q��C]j�n����G]��}�W�tϴ�T99@�)L�EQusGbV��:\?z�8w[����x�6���wG�vu�kQ����n,B���}�6/��Ҩ;2Ӹ�Yn\4���D9IÔV3�lp�o������P��rw?�#
�&�� C|��:�\c P���0Εc\Tϒ3�o��ʗw��u�W����X��{�C�z'������:�'��W1�Ig����E�6�)+�DG�n��p��Y�R�]�P�1�k�3<��	�qD��`�C�\�G�E�oc�D{�v����[���S2@��3ڻ����5	�$�gB�~%��{{����|eC�i QY���_��)�/��3�+��ȗ����8Wۏ��6�d�'Ų�n������{���gAF°,q'�p0oܬ��▃J��oi�_=��M�p�։a����Ihj�(��0k�*	c �5tP��ݹ D
懆}� ��N~���9#P�)#?Î�*Oy%U�c��r<!c��ފs���*����@�Ɂ�r�L\q|&5���r%���$],��6��!���b�W`S!l��6�Ӧ�e�Bۑ�<[R�Q?���66q7:�s�n�����P"�	�Mr��Q��t�'C2}_�;۪Rx��S�:��}�!H�ւ�T���o�C�7/�-㐒�ǟ�బNA��I52��|�5ʈ�ܳ��%��I�kkG&���(��.����MƱ�1�i,P��㙄���_#t�!�>�$<|w�\�N ��2A�/�>5��C�A����F�8F��)̞���C��bj��Q�'-����?�a��?����7�;�]U]%��	�c�c��Tt����&q> '^��7����������ڻ`�}�/�ܐ�7ײӣ8f^�{N�̘� |���� -b��|�3�r[�*qj8�Ѧ�s$��s�u;T� 8Ę?�_�0��/ٯ���s��`�ӣi�ӑ��#-	C��t�Ȥ���C'���G6:(�p�˞߯���}7��-q">+�
��5
I�A��
�$�1��x�ǽH�4e�G���bV��V�>M�H ����Ǉ�Lnјd Pxm�|(�r� c�mő5�U�2i������P���tg�ne~TP�}�6�^�N�{|���9*�g-�\�F��6��[�9c/|=����DXDB��	GX�J��r�����#"���q��=���6lo�Gj�H{�b�y��RX�mi �`Y_&0k?
���7WGG5��F�g!H�L�D�'#5
���'�II��Co���L��ç��0?!��.ݺ��|Y�c��!�<b�5�BX\:�H��,7l�