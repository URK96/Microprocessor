XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K�<�̓l�ܔ�ۄ��O{��S�sЊ���<WX~�����0S&���E�����:<{�qC<w����t.�LdU�۴Wf�^i��܉�a�3�H�\&��YDmI�� ����u�I2�?7~�1���0C*����/_ڻ��X�N�%���	w[KJ�x�nr"�cs��b�ɻs_wN�m|�۝���#��)�Q�A�yq�Aٓ��ٹ�R�v�-�B�/�&�;��c�K	�['��ͅ[���aG��O�O��63k�3�t�L»�)��LDhw�kU��!!%W=[ǹ�Gf�"~4�'e?W�����`�;.O.�A>bh��.C*�3L���Z�.}kQ���4�5����/�e��
W8�����H�"@�DE`+�45N�y+�؝�\o2�Te�~�3����h�M�z���*~���{˦��.HVi�������P'J��o�w^WA7�G�Lw�(�� �n�EA����E���=�-}{q�Q��Ɔ��{���7g��#h�B�l��Wj6A���w*f���W���HR�$?U��H�:{oи4��� ��O�- �;�i��S��|�99z��F8�J�s.�k�hSz�Q�G��p(h5��-��ɳmN�`Q��s�ξS:�w��O>�	��u�ĺ�L@�.=4��ľ�2>�ˁ��������i�� _x �!�jȣ���Ɠn��u�F�������T��I�,{��NM�4��]�O�R8d�^����������
1xcDjo��A��?��0^�ޞXlxVHYEB    3a1b     d40���X+Om�$#��"�H�M���9��71E�}�X��x]�g�ʐG�Q�fLb�(���������铩�kǀu�˷ƢC�7dKa�z$��Q��,4T��s���g�ai���=�X?c3tx�Ot.^.���'wF��E+~}1�g�������eb��b�c���*m��� z�!�|�J}aV��~��i��@��c�������D���F������Y�=(���J��(�Q�D����͍Jʩ��V��*�4��������:�ʯ�g���,�U��Gq"}�E�����ܽ8�s����H������R��s�ݓ��"ӻ�����������e���X~�&��YZ���{g߭�.>�fxL�yd,����2|�R����4��.y`��w�ʖs�m$�3��T��T�6+�ҧ����h� �nmʂ2�As3JQ� Qp���b��dRP3���DU�5mK�MQ���V���Uӕ�+��6�1Q(�>�)Bs����4R�_�Ϸ�h!�=l�xM�񍽝��6X���d�j%�&Ö��G����/ �Գ���Bၴ~�&��`L��d��g�� �ݮ�����<6s���ȿ�H��*��xT��!�]���<Ϝ�xk2�۔h/����CZ����9�-��#����z4�.����i~�����aw��8Ł������
fe��}:�/����~j�����X�.rGJ�7r�ؿ�ǖR��D9�
?���0��Q�F����A�8h��x5��NF@�FM�8��-)b��?�������K��z%h��zt���e���T~�gk��{C�{�(���e����;JQ.�� ���T�z������3t:X��4� �7�4b�����<CZ;J\˟��g�������m�A���V��h\��һ��S}P��[b8jp�Y����2ƥ���\��^/t��/�FE�%��́�x��S�̲Y�9qQ-m�����Jt;�K��7��g�7�<��?�z����(&�[dn/�}Z��b�b��a狐ѹ�I�LO%�c�⾳1��t�o�EE'��J��gvA��k}��.��Z4l3��}���1z6�r<:hJ���������4~2RY���倲�\&�o�Ӟ�4z�sD��X4͛�v>,>����N	��&�����!�2c(�T�8@�&�yH.&<�~Ւ�`q����x�k�b�䫄Vj�����H��a�46џ[�n��2�U��ZB�c�S^��7H9A�`9(�����7��Lzd�$���h˯Wi��rX������%�
�#cn��Fw������ܤ�K�A!��:�����	7�j�|jP��\
�6(1����e/����	G�{��I�K{�˵�����P���ܶʋ�j�X9,��6�[�K���!c�iH�����oy�K. E���겜��v�Ci�&�k��Y7��E~���dv��O�D�C}����4�8�s{2cF�ǽ�6�W4 �U;�w�'*�0�����xw��m�X>�����5���6���j��[�MI�}'ɳX\5�
L�p�=���� \2;&^�� X"4�a�[a��3U������?V��<�5dW�/
����d~����3CA������%*h�s���q���a�B�"46Z���&4�u\&�w��w�Bt$���EI	���	UUJ�H_��4����Y��J0�AD�/}x(EŮ�+�G�֒1��/�����P"���.���5�s%�cv�6$l�+�>X���@�h?#��yX��tQ�eA4��lC��Pt��
��-~Et�o�D�L�Tt{��4�ǻ� nb���6�,����,�.e&Qi�|0���:� ��㏚?9�z��������7	ƙ�R�
��=�ؗ8�sVC�(�eXLę��b���$�"H�N=v����ܥ��$�K���!C��db���,����֗���Ib9m��
�O{� Ȃ� C6}�X�ʻx���ԫ���V�@I����&��@�Y�C�@7���b�#g2eM��^��l��T/"������3)փ)\l����>�'mj���z!6�BkЂ�(C��7�x�:���pt�+���p{��`4r����s�+/u^�h��S�%�Y��PL]c����ނ�,N���^U� �S� "B�+�Y��C��u�Q������>��U��o*�{.A�0�'F(F��8��A�~UfL��^2eS�!uM�KPD+�g�'�n/��S�5M95���E���e6��L+- 1��=q�@���z#��w¼�@.KC܌7��󸈪�YE�w�UV�5��L��A��?˱,��G5�O�0�O�Z�V���s=$��Aj�%�;Т�Ɨ-���{N������$��1ud�a����8���V���5���x��a�HEr��pe	�~�6ot>fH4O��L�v�3$�c䠀���,G�Yk�!vD�Y�(�͍�g-�̅��KTG��U�� =b���I"",N�<|�l`y�q�j3�*�Q���O�E���CrP�E�`
=��G��'�����6�X�����F�I�2� uF��#x�p�q�����<�65���s����/�a�"�2�y��w�y5�DF�]2Z�0� DR��d�&��p��6��&`�<
���'������Ȩ�����Q�kS�@�ܩ1��\Â��<a�a2����8�G�L��6 ��Y�����8�\2�7͔��ϛס�j�]X���*Ɏ�������=��"�����W]u�E���`Na���l,m��;�#�c�g�؂�9�$ �kS9V�-n:��.�$Jɰ�s�?�@� �W0G8�0������q9ǜ��@�]jnۓ��?�X��QJ=�g�g36\p{��C��8%��$���q���䄾���:�eyT�Dܲ�L�4���nK1,�y�B��c)Z��_F;��eyH+]��f6	�A��`�]s}�r�S5�uS���G��DΛƳ�E�F�f�wg,P_�ρp!
��n�VF�6B�\�$HS�����[�*0�_�[���xպ�o1?i��DI��r��B���� H���S�D������#>�K#)mĻ)�|,��fV�{q�%ޑ���|ǋ";塯� ��
lH^��]5�2 /:�Dp�ң0���8>���bdE4J�&�T
x�1e��Cb��ٟ�w��E��ד�Y��"5�t�6�J�+3��9֖&�f��]��|"�m{�n�����g[�B�m�R=�D�˹����]e�����E��3K�ݺ�V��b�eQ�kp���<	����V�����3Q����β3����5��Y��5