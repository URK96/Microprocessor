XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���/,U�}�@�:��K�oa�.��l�Kc ��ϱ����.,��������&���F��|,9��CO�j��:� �Y�#�y&��3�.v�z�v��GQ�!���QJb��4�D'eյ�����ʞ��$yK�'�ۆ\��_� e\��M�EʤLZ4n�'��sY�m��4�
�^K���cHw��&ߟ!����k:�TcM_�	ϾQVNK�+�����#�EJ�$;�"�Ɵ<��,��Td��nU��:<�E�_ V�T4/W�3���.x�Mи�TlC�].�&�',&��a��B,@��>u�ǹ���{H�jbH^�;���M������ �������Eк��E�X@VE�ň�q^p�IӐL�}~Jd�ϛ���?�kt7���%��s~<|a9얐�nt�z:0�z�
Q��+�2-.��Ղ�Q�O�ڌ��	Xv���Xx���W�jni���Zlse&�H��F���֩����[�>VX��#�˄Hn�ۃ��H��J�&���z��%�ڱ�JTF��, �&�tװ��� hϣ���>�@��8!':)��*�&�L���]5#�UyW��=�6p����ʂ����V8YQj��4��P�~l�n,��b�*��N�Y�d��d,���-=���5�!�ˋ{I�� ��
_ܻUo"�w!h\�B�0Tԧ1�±rJ}������\�Ju' kP���$�`/���ɟ�FyHT�L1���&�iy/��.8�e�zh&O�4h��ł�<�XlxVHYEB    4a09     920�f<B=ڍö��:��@�[�@f�4ʂ�a���r.~��!xan�l5��i⹯�'�k/f�0ݛ���1�u��W��σ���V�ڌ���N�H�[�vu�}жl��/(����1�u�j�#��-&R�1���j�u㒠�8�.�ʉ������mZy3<���	�aCwK��i1<z�~Kq6��
���Xz��Y�Bʵ}��	OJC���xf��~�OL�u��t6��
Q�-Vޔql� �����a���:���uӘxY
��:Z'?b;K�JO( ŧ��p~su�T5qL��l�$�^�~к�-�k�)ǆ���A��#���wSb����/�0�q�QQ���f�s�crO��1�Ī�9ؒQ�Z-��T�W*�ZqH��쳃O�g�F��Z�gR��R��1;K���N��j�p�O��_�ӹh!����S���*�t��6�� V廙�_�A��㹛F�"���� �`�T]E�^9Q��,~�s`+�\�!
B���CF�
�o��3^b�Ӂ�Ć�r��qH�B�'� �g3�9��h�()[$E�`��&q і7�Rr���ڻ�N�}p�LQ;���8Y��K[��T�EKh�*���r�t��f��5=?x<������Y!��˕��X�T����%��=6g�.�Y��9�)�KP�J\�hRǥ�\��ҸU�GƠW5�?�E��nӤB=���!�^�|��{X��>(&�F����>>�����/~�v��#:�@-����B4�q��r1e�{��T�2+(^�0P��;,m���v��G�Y�zF_�3g�3+זe���Dҁ)��?�>�q��
�u����eei��ز��r�ԧ����/z�N�����=f�.����,�(�0эq�8�L��]긋�[ցh�H��H�{���yx��@�:���^�C.�+C0����u��3GX
�9y�߯�Bo2�Ӑh��Ӯ_�Љ�Wu�߆�\��;�)��5�fjQ�~�B��l�F��n�Dh�w��:B����ά��-4x,-V#�1P�O~��?��g�o����]r�Z��7s,�:ff �
�wi�Z�7%��� :1F�Rb�&=���!X� v�9A@YQ�%�E��x�rk�@;�5yG��L8U����6(�R��6�D~�<�,S6} �CP^9��L��{#�������-:;��ڐx�}<T�lj��5UDV��J�]N��H��i�y֊��l�?k�i�ؕ邦�Z���.a���	u��5�|�b���20���(>��!dTB!v��^NET��]=�	D-�ؐ��7�c��cmʅ$�F�����|����)q4��jP7Z���C	�L4ɳ���6��E�4�������~_E�j��GI�˰�`z���!S���Z-�K'�+�}BG�8��o�N��)�	���3�ؙ^�-��y�w�piwE�Hsk���;�f)6�8��ܾ�P�Ok-���T�����?�eyG1�K�Zk�٢�3	�&kJ�k��m��;�p�R�a#ZnYP@�&{�n�Ȋ	[	,-���Y^�O�65M��YK#���,��I��UJ6E�"�a�p	��<�Y�
��Y~�U(�'f��� �J��b%�M�+�(RJ#)KaȬ�a�>����ͤg�	��ZS'�<v��pq"?�{��;�%��GY-%��H��q�zFp�Anz9�X�]��&���TF}e��qi��H�}�0l.[	`��Y����P
0����.��u	�K���X#	�"�76l�t����Ci\ [���ú��v<�W��o��>��(��LJ�OЩ��_>��X���ɱ�.p?R�j����ڝ�*~�
�����!u����8Q����T�Tڃ\#�� �k���koEiz�Io1h#�$Dﮞ-oy���!(��I�+:Q�n�@\�{�c[����7g��cuM>6Ӳ큛��_��x�����oh���,5�������n�,v��!4�����i�b��9r��w
h�^-�ʼ4�j���"o�_d4Dt�%�OvY3��}0k��z7�T�L ��.�����Đ_���R6T���u >N\� 3WU�/?pio�R�����]��]����c9��PK鵘8u����A�&�_�m�;,'�ש�$����=��c;�Х��-6���l�B��|W�J��"��(ݺu�%C�~z��p~�s���fx(x�|[�}S����ƙY��'Q����v�%f�v��/���s��l���A%rn�� !9riT�S0o��pp\uU��t�A���-a&��Ӗ�g:��c�j�����@