XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��O_u�^x�W�^�gU��]�v쉖3�����S�Q�{ܴ����>�y1G� ! �Q���5Q�.J*��.��ge��4�g�V��P�.bE��&V<wg�/û!�C�`i5�b����k�ԘN�Pj�Q�Is�K(cՃE�	�V���c��ܧ�L"%$�T���N�1FxW4�ӎ���q�bn��# ۗ�@�{���oK�E�񢬋)����]��q.���Ś�߰|�E�7A�Xʤ4=گ�&��E��a��L���l���6cs���f�`�J�yidx��K���C�����}�r�8>:+
�8��Łz6�����w�]���$�	7IF��͢~��R@�xN@�r�/ާ��0�(�����9��PG7 �pc�>��.������2�=�8���3]�x�,�����qD%Ogӳ�I�pU�L���30Oy}m�V�HU��Yݍޚ;��l'G���g���VzGi��@{Tߙ� L���4�Z8<���Ң��p�IC�F�g_�/�����"�6�L���cʸ�|���� ��8���v�]��`g�m�>	��$��OE~oCr X��egFqE�*-��̩���a�d�o�ZO.�'i73�����Z�,L��L��D�N�j�����TUt��$14�*.;e�x ���YG(�K7����a.y>��܃�*<����XH�ܹлy��e>�jZ������:l�������� :+v�������g?����O�+��iE�"��>i޾bXlxVHYEB    2861     8d0Qr(i���KvE�pu��$��=9��h���Œ��۹/�������+a��Q>����� �Y�t;S[*!<b �����U�Zyp����O�~�~�"�j��G����&�\���z��G��-����&^���7������ï��`��4�>#M����L�4)�����g���ZYM��]�{h�݌�2�2�%C���&�~���:�����+g{�(|Gz����k�%�|tҬ���_�.7Th\M]�F��H�' `�#x�T6�`�qLݤݳ�n�֥��F���= *&f����x7��\Ɨ�}�BБ�>D֢����x����%Sd)q��_D��6���؜�� ��=��T�_0��?���H�Z�/( �S9�<��8Xv�����H�U�[x���47_D������8A��!$�t�F��[;�,�>�}|f��yk-��})m�B7��T ~7%�`�v�)��8[��Qp!3�C�ڂ���_�����$c�	c#%P����m6�s�Ix�dX�u`?�W���M�u?��.L����|�1�G��ƈ�2��>�#��7�Ȅj�)��@&� f��rȗ�g��Q��?����	�E9�eT䗽X��)r�8�|�F��|8!*V��t�!A��%rak�C�Г2�*❮��ר�魋�*���������o�+��!aP[a��Lm�5>�#l�����"�:3���[�0Xݏ�6a�n}�[J��	�5��*�c�y�Ui�I]L5�[�(�t����|�����#ۇ&=�-�:KA2Xn'}�,fLH����~�("x�j�$�����KN�&�L�xU�B�bk�A=��ly-]������?
�o�7b@X��oSHP�ڿH�f,� ˝3�/ �Tc�ɐtgtuA��嗷��]��D}j)�$j��ʣۖQS)�#���Z���o���\��-C��l_`sz�S�����MhU�EmEψ�!ȃ:ۣ� ��|�������A�E�j�����mS�c-�U���B���@���%���=�B�fe�[�)���:q?C̿�ح�WF�)<Y"XSO�PK�K>C[��h�����Od��'1\[�;�|B�ø~Q�J��[��Q�����`�܉�D��� �307��_��Ͻ�v��V����;��}_�E����%D�DK�:҅Mз��|��T�i�!08g�^�a��l3&X�c�Hʗ~@�Q~@<�������Iq#�=�c1��6/�6� qtr_P��c��e
��g\�UO����JN��)F�b����#oؔ>�+C���r!xPb������68M>=��6�lM�����T�p�;�]�9C�����r����å�+����Yj�M��6�bS�)�*a���L�:;1	ю%gJB�/�]v[��(s�K��B�T+qѸֳ�ա�uAiPN[�!9K�J�->�E�����G���vWP �Su�����A_d$�4�	Î%*��P��D@�f� �H�sk�>%�D�(񒁐��b�@�K�~�8�����(���eI�)3ɸh��<��}�k��W1��Q/j{�����T�@���ĸg��'�F�(AgI���]*y�^,ҨE6'�ր�L)��o��zNMEŉ�����װ�u���X��Oos�hp#g�KȺP~�28�Z��"vX��<>7���tO��#�s�O��Yb�t�����X0���w�E�z���&k��t��;��6Z#�^m=ݼ�0����w��`T�$r����FZDsYJ�;f�T��H[R],0��0��ù��kLB���,�<��X�R�K�aܦm&�2�?�RX�� ��xˍ��Y2��b+�Ւ�σ��y���N�x��P�4��'/����@����A�Q0QP�tGn�Bm�4�#�� "JW��K��Y2s���t�K8b+Q5�g&�
�]��7��q�$��<@���r2���!�9�ͩ��)]���w(���'��ý��V�pZu.��h}�e��ʑ�5��\R[�>���Z���o:1C B#�L��,��F��W5�����YJh2��ϼ��H��.n>�wlW=��O3���uϞ�Y9b5�)<�7���9?��-�֋Э ^-�`���S�N}�'"68N�s#��bK'
_9�H^�F5BK������&����0�f��B�*�y)��x�8�^�ƛ��<U�x�
6�A)q�P�B���(=�!�m����}Q�X�|���>�O�&~��{@C�fV���