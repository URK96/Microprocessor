XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��qz��zQw��=�g��<�zw�,�s%�D�_�~��0
����{�R��tv}�: ^KvArS���5�N�^f��I�9F��pajΚ���4��;�MN���R��n�H����􈛂�8u���D�"K,:�p��쑭����I��$}� ω(���Ǚ%%1�����)�\���{l9�W��X4B�#V7�� ��Ә����5��P}P-�Zl���!^��z�g��6�r��Ȭ��ܞ�zuS�0����Z&q2{T��:�-0��w����0����x*������/�l4���th.��m��̙Md��S�\N����r �`�|Bs�����^��}j(M7-�E�u/�B���=.�X4	 0A�8�㠀/Bi����3ynd��@�\T�{+u������2�$� J�c{(��M������n�`�N�$�����װ��.;4��Һ��cwLU�'���4��φȂi^bp��o�C�Zio�622�{���I�*u�lc���|K�qzל����ᓨ(O�4է�-�\��-p��K�_Gφ�^���gm��/AS{�48��[����
��	�߲�������';! .XhO���RK�
�P�2]?����Ÿ�s����L6/f��:|�A?��;n��Ɠ��y�>��4
B�b)�@�D-/U��}y(U�%)�1|�v�3�G��5S��(�!*6<>R�K��\���*�Q�Y�G�m��0u���\������6ԓ'PdxH���\"��cXlxVHYEB    4e25     d70���'�k����zM����_��c��y�N���QH�-O�'{��-�	f����he�w�%�{e�f�pV��6��検�zy���
u��!�4H�6i�S�Po�������[c��h� ]�����=�+hCz�Ʀɼ롁S���,�I���i���Rc;$%@��3:��t���l�����e̎��� ?��s�7*?sck�ö�u�m)�~y�AԬiMq�[a1Z�>f�k��D+�7��=- 6�c��� ���O�1A��5���h��=�g��V��
��A� J�hi`7bs�8<��M�W$Wq���$�RX��wIa��^0�y��IW�Q@	(Mݮ�kPs��m��I���)�IWr��rT+<�r�)@Rx2c���:#�����\���il�du:��E�2W!�c]��ؔ�XT�~.f�m"V��u��K^���+V���fh��߸�v�t���XɏR����#]�r+�qv����KvB���,N���A�D�s��i�!���i�5���
Z��~�`k�&����ݟE�DC9�I�ZS�j�����r����&�V��4g�L���Q��h��d�FTۮؗp��'2>��x�x�X�|(A��a��ӂ�ȴ�S�sa}�G2�� i��Idcw �*�-�R�?<vL����Wt�Í�h�tfYUAOq�8 ��󘓪��.� �M�Ͱ"��vQ
�%���ص�޲=�V_&w,@;$�2S�Q���l�Y��^�b��5�m��d G�L:�[6�H�e����5"������jhe3N��?C�]G)0�B�N����c�0�(�*�'D�6����>Tz/�Q��W��<��Uv�Ԏ�^?�U(��p��8�J�P��Y�e�*e���]��e��q��0����Y\����|����z�.7r/��y��f����`�5�oVU�:ɿ^Jɦ���_W�z�t"ļ|�R��R� g��n4�)��������nK2^��˥T���՝�r$N	Ւ�F&;�t��/��[��ȝfN�#G�<�u���vJŻ��	yq��r	���vh!�����6�Za*ݫ�k��sNb�%���!�F��wc��� n���\`l�!\�ɋ���g�V����f&�i�k\�Z�E���H�&^��#��s��%��:�C	
�7#X��T� 	��Ip �@�g;�&��n�v�O��-�Mp|8^���2HD
�k���9.�tZ�|��mxy�jOl�~tE9)Zm�[�0P���#��UU^�5pdr OŇ���e�cc�r���'��/�7I��{\_��q�mT06�З8�1^��H� �p~��?^p �����gUM�ҩ�_Qd��C� ��JN�*�h�_C��W�eg�TX��z#G�C�>K��p��
�^q	g
4�=sX;i��9l#A'��5�{'�Ϛ��\A��� L$o���gB>�$(<�y�%T@��ca��υ(L���n"��8���T}��Y�ߑ�v�x�<�3A���wO��eMN.DR.���"P��"k��3v�mm<K_��+H����rX�Ԓ�΍�4.�	~�n��;���Oc,y��|O���i�uas!�7��̭}L�4��U�a��k��F��+k��������j���H-j�O� �����p�5S�����̅x��h���8�^���dEJ5Ά��00uU9n�"�nR����U���s#��e?�~�A�t�lz��W���~�)�$��Pi�촣s�~l%z BG�<_��mH,�\o׭=K���!y�`ķ������F��vNJ`h$����"b���[ ���f��<��XPr^2�.�5���h�H�0I_�fRSv��������qJ��Q�Q��]&��"a��u֯�U
�=����%����킹�g�N�u�Q��R�oV��/�|�Ku�E?t�w�8�$�C@D͘h&[�&J�(�8����I�� ȓ�̔jg�r>i|��1���L�@�/m��f[7�A���2#ݡe�F9�?���!�	�^Kj�h"��������5xзV�4b��w[�)Lc��s$��js��&ٗR���)�D�D G=D�@��SC����f���}]8?�:cd��?�t��l(�X�
0���l-�\�zTP��dM��mY 0��4_�'\V1,��cdE��r�0���|��
�AU͸_-V��5z��E	�֌��l9&�oN���y����تk�Q]�i�Ίۭ
u l���n+O�L�5JAb�!�tߔ��m�&���ѱ��U���;���<��>���s���y���d��]e�s��@Iu�+����x�p��:^�|�:��R250߷�%�ՠ�h�z�Ȑ#��>G+��_ɇ��7�ԫ���l�`Jь�z�f;�Jק3�0��Y��y���}˙�+�9�T��gץYH�#��m y�IB����#{����Z�e��U[:l�c^����y��o�D�
�u'1c���WA$|��Su���l�d;�AID3# 1�%�+�)���g�p0���Y�/�9�����cf`}m_c��7���[��o�{�՜zw<пU4X�TyR'wߔc�l\�`�h�d���|�lf�3A��Z�C}>�ż ��Q9��ꈕL5jX��eO�:�4�B'Mtb�D���7g��)V�AԘN�_��z����T���u�3��Q��_�=���3�?�^X��� o�_�Ӆ��}�|@�\j�N��F�lY�>�P62c��
�-� ��إo��1�r3�7�ƞfW<̮$YD)Q���Qg��v������X|��*�}Ar/�v�N�wJ8���kl�4M�����K�E���Ͳ�-�6u��O��B�c�ͮ _[pu�gѺP[�а0�ހ�Rח�0#��"��x��� �7{-�Z�j(ǜ\ɍ�ȏ3�۱?�yK���
��p�J ���u�[�V���DvQ�h�UE�0����q�[ 8�U�k�O�[��ٿ�+�6��2-���
l+1�i����Ap,���[JRU�	B�4�q�p��Gn�$�@"=\ �mj᧛9�x���8��UZ��zɪ8^�W�40�
����Xz��D|)P�H�d���[}��æN����^Q���~��p��bK9�ʃ�(�|^��W�_�],:��Sq@��u��䅬�IZ��q/a���69��Z��*�b[x�Qۖ	�2A�����6���� ��%᪤�>a;|*X!��v�^j^<�h2�.wa�6�TQ���c{��)X��)ڝ��l�ξx���{ �mdtVR]�B&bV�Ƽ\�sa��«��%�t��-�azo�등����Z�ހB�H��:o��>83H�2|�]��M[(�(RS@>NiR�́