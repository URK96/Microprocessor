XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���٫p���#��:��dp��K���7چ�����O����^(X N�����):��7��a�V���� �Ȍt�i��-��* dN���@��
D3[�̠��8}�3�W�G��y��*do��c/ͧ����6?Qt��!�:�6t��3��xH�T��U�t��t�d��z��_���� �0!áQ�m&��ͬg9CS�:e�Z�	m�n���ߵ+�g4�L�B;J�a�^�
�v'(�6Wv�_V���;��jh����/����7��]
�+[�X�{�G��c�� ����z��{��Yy���M��:����"gğ۷7^�g�QN��M�l�-��o���X�g8�`��U�d�O;`z;d־ �lm=}�@DM)NiVߜ�@��D}x[ǳ�P�:��B��T���}7�`�����t��P��`_�ݖ�k�pE�%`�Hԁc��dYPa �9�5���{��|s���Pl���D�^)v���9h�s�e�_�c�6��,�bm�9�:L�XWX�s��3���6�Ȇ��ޫ��'_}Q!�F\�|1,��C��
uԸ�$�����/)x�6�$dX���b�mԦⒺ���3s!d�1Kc̸��S*X֨s�fs���e�k��}aߌ�5��(�޸!�x�S�%�~���t
�
�Ռl-sP
�ж5#C��i�S�[���Y&�|��;���pO6�vo�e	ĩMH��xc��2�B�]�\I������Ρ=z踁$U}�K���=>-r3 �;X�XlxVHYEB    3246     990n%�
2�cN�������� N�j��\G ueY┷9o%�AOҽTiμ��P�����,߻�`�W(U��q�8�iF= �f߂2�o���-��[��GDc��&�\�LQt*�:�������h�=[qS���TN@)ٮ�Aku" ڕϪ� �j�6F�~��Ѭ�Y�w_Hi�6�y�jO�T�\�W�6w-��ʱ�<"Z�7-�ك����A�4��m�-Y�;njm�p�(�c]��S�/��,�����I���b���
8aY�L��-
�vJ�������5v_J祑�g�¾"���fؾ�H4SU�W�=�0��0�D���J��kt۱`99�t�ƛF��2 W��ϕ��G�E|"7O�w���eV�#)��q�چɴa��yJ� �Ңc�J��^7}:�Y��(����#�+^�����f�c�/ߴ�z_/��@}5=���G4�f3qE����B�\�v��"�'�՛bw>�.�}����i�V�\Wِ��X�H�;IGO�����6ԇ���Ҭl�E��wx�h_k�yJ��>"H� �Q���D��s祖���0��&(����qK��V�1.��a���x-�}�y�"DM<���b�1�Z�v�L���m�;[��e�������h :K��U�"�OPل�bŧ��!Ɣ�z��0���<�ŃҘ��n(�89��'I���K/"t�1r��"���&�u%ocWl��_�5n�UȨ�͙Rnt�t�����v��I��XA@��^4�;XS�p��	����7ÞC^ ϭ't l�(� �3�Y���!y.��R!����낉W��(՜���������-��+�>SGo��H7�͊$k��%�bi�� �A����Ψ[mʥ�y�zOJR����ǀ���氧��T%�����F�#o�̠�
�Ҟ��yQ)�"��a�?�4�v�f��-o;Da�7��쌞����ͩctl2�	g�2`�S"k:�o�#-T�*ԧv�Y*f���y�"aK.��z�;&A�\J����>�fL��@涯��_
i
|�g��~�_��V+b���{���Da5�U�[ֳ1��w��L��$�KB�*f����@#�8uʣ.y�M��H���u�EP.yM%k�4����vH�pHg�E�����ƍT�7+�sΑ���xd^��T�#�nvX�9(���{S�%Ή\�� S��N�W����\ǫ��-u���;�%�����*���m�}�
���LU`bK���sȆ�e�<�E!��v�/RSNͧ��*Wp�4����x�C�^�d�(�4��m����_&��(کE�
��V&�	7����U&�+�ed4��U����ވ
F�do~�<�5-k^(Y5��,��,�����BƳq ����-.ތ�?B�X��߽���B��Yi�&���7���48��������*c�U���a�@���ecTMHϦ|z�9n��x���k3��@0�f{:ǘ�_�*�
ρo�	��,*�87#-G�[%б�$�w�:��3g�x��r��x.}�D�R��q�+��[ ���xmK�ij¬	u�19�$:�+er.h@}�m�r�g<H�"�6�2x/~��n۲�D��A=�W�vZ���qZ�͹{_B��v������'�=κq�l �v�yp�9O��M�!����� ������J�ku�$W�GK/Nܝ�{�
��z?G�~��V��&m"��?�7�g���z��_j�&	(-�B�\��(�5��-}Ծ\����_�R���hR��j�j�A��%Ż�Fz�y�zMŲ���^?6���{�T��,w[,v���)�o�Q��2�6�[�
q���ϠUNj��0�+(䎭��H�"��e�]�Ƚ2��g��z��g��I���I���q6t���]�q�XC���Qf���_}Kwݪ�X\����aW���d��^-�[��+�|V��>]��K[��h�@���4?'M�E��A!f<�W�yV����Mi����[��@��Ξ��ffĦwo�s�VZ�����U�T����=~}�b��t���E��P��̶t����)�U|��>�����%V�$ãW�s}�l�d�5h<���7��4�f��]���Q�L���I�|��egS�� �3���l�����p}ScE�T�J���͒����:��
UrsH�cq-?0uZ�~8�,�d��T1�Fdщ.�kmk��*u+.�h�lB�	v��T�Uɓ��\Rd�XFg� U�N�a������|+�~J��d�TW�%�]�a�$��?�%E�@��U�P)�y�<�b�E\n.*���rM���_-�<��h��/����� ��|�>rZh�_����-�C�%t1 3���ol+#�q���%��iz�Vl�肻��(��0׻