XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���<�z+ ļk�$��n���(�E^,��B������_����:�!�W�m\��8rv�d!�������|�p�����{@;�������Br?�j�` ��-Um�����2�q꘍��=j�wd) RR��%]�1Q�M���M<��ǂ�i�w��~Z��q��zLә�)�(m [�F(Lߡ����m�)V���8�Gt�I'�"|HhF.��k	)�R��#uS����o���e���GO��Y6;�Dy�� �~-����"�CY#|)�&{j�\�FB�s�f��	��7*���bz�k�{� �A"��4��.fM���V�߯[rI\�p���]�ɲɼ�s�Ɔ�K�R`.����F3,�-s�O�m$ҡp�x��#4Dl�=V�p��X�9q��3�G�}y�l>�T�a�{��n��<�/�V�vp��5���M��6�����29kw�V�)9�#��[u�UE ��6�1D�.HeX�X��,�I�x�!��iy'�=�ܜz�җ����ޗ�`v�n^��o�u6~���X7(�pW���K�4p�V��UŠ��E��UI�MĀ2�pS�<c3��"|*�8rG�(4��4����4۵e�O�ν���B}[@N�k	�N�8�T�|]53�p�l��fڱ�:�":�:�v�d��u��4��u��?/�p��B��F��6
����'��ό0��`7��M�8�*�u���Y3�#"�������mX��x�u�Y��2��p�XPk��
����F����mXlxVHYEB    156c     590��=��9�5q@�>����D�җg���D<�0����T/-N���pw�r�)�:YT����9,���-d�	����T� �&��{s���W�e�z:���wG��W�]rd�a�83����i,��G�Q]?cI�N�w�!��S����]K�<=�x�uMe&L��XN�})����U���z�'x�O�i�E/��|y�=�[��wXN7�k���F�A�i��L=��t�9����T�T�'�.5�yA�|�oCmL��L@����k5�Θ�����H�7 ������u�Pc����<�G֒�5C�d��ʾ�r֠���,���\�<��xVe;j��O��ݺP�s���4_�?+�O�T�	�6E��闣Nm�m����W<�����x5��^o"HR��.�R���O¤.)eBi@�(v�/�j#T�Y,�y�Z!n��m$h��g䘙w���}�j��ŧl�8- �s��]8���^Ri�땍��;���X�������_<�4���ҺX�%��&%��Dp�W#�T���h2��=�~f���kgJ�M�y-�!��l<��)�2��S,T�	,��Ԏ��}��bMJ?f��o9�V(�s�5�kا�iz�
g�Y=-)�@ۅܔ�'eR��b'��|��N�T*��%q#?�.���Gī%��@c��2���������}�Gfn�����&�9aYݛ��s��tU���Ƒ�!L��D�"�ᤨ*c)�P�?g��m�^�����a�n|T,�����X��ѱ��a%��T�~�R^bk}[:�����+�/�Q>�[�bD�=WZa�LrB'o#�j⟀�*�ao�%�+�:�㴼�e����J*xP�C�������*в�#{8R��\=��uUW>�[k��.t�x��F��!���T�
�_@��'����ay�ß��m/�Y�������3()u����[*~�r:&�Ѳ�V/�~�"k����}�'F[11=s�t[)��fH�A�O>"��g��������Y��/�2B�!�w�d���z�N[����Eky8�9������q{��T��zPW�_��y���l$a�o -xOlN��U��w)3͑Zla��s1"Lq���;`���/.ZT���
�QM��X�-�P6�=H�&�5�c|Q쫻�y�F��	H��t�-��1�?�${f!B���P\�@���.�l�ʱ��d�=��CU6����]T�w`�B{����T��&8)����|���R��R��,�TF���wd�b0�J}$��SA���a��K�FT&�<f9�j��%K4�[ަ1=5¨E���u}&ƞ=h��nu?���v ���OF�_���Ya�����G�p��@�FQ��j���6`).