XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ika+k�-�p[�~<X̢??��ފP��(�M�сsd�n'�0�(p��=q&���l' K���� �~��x� �{����Ai��d><ځ��lA��%���3�����js���(���穗̨�qՑ�	`Ľ�=*[Y���@��Y�Ɂ���� O�#+�"f��`2yGXT����A(��K��;�V���G�0p��G/�[���hz2׽'	/H>�^�@z���2LX�������J��Ţ�5H�jb'9&=��y��)�-�������ءv�Ը�p�kp��SgC�ۯӠ���85�\Z�����:��'�Ŀ�͉�(��`�T�&���럸1�2gnK�T]��w���Q�#K3-zo���j/�o��1	����:���Z��X�w��qx�m�*�z�J�l4�r�j�4\'�����:s�d�٠.Aly�O��HsG���x���I��qq>-&�y���Y�Kgw��.� �UhFm�G����'�2ܽ�J�m�U2D�&�!��'8��V�%�F�S�n�z�$G�.u�#Y�}�G8���\�F g����f.2W8�_
,�Kػ�'h�S��/��9#=��1؋ҧWF�K1��c�?�^o�����5!�ke�%���<��E��i������ua�=�)QE�+/�H�S���U�[�����I��(��r����/���@?Tw9+�=��?�,�<���h�9/"B�YF��Zq����2���:*&ڰwI\�6<�4_��k�/G�(}/x�����7O:��XlxVHYEB    152e     5808�y���L<�-zС��<g�.�F�8��g��`?�,E%o���n�]�5�ڎ�.�E��vd,�k�:�6�I9�Y�Ȯ��vC�0�cʪ��E_�,���_40AjWG-��Oh��{�IҼ�ѿ���c�H�
�+�Q��B%D"	��8Rx�c� l�l�_����L���C�A���1�#�(���6�R�8�M#��� ��Y�W��6�_��SD-Rb��z��O��=�#�&���A�]n�Xò��)G|M@�KQ*�΍w�N�Y��٢��sW����lW)Թo�^�@�=.���s�\k笜U˪ِ2����ͫ/����p*Dڦ�K�Jf��Da"8�wE��'�V D@ax7�j~�W���A(��!�o��mL�k�*Ck�{x9n�r�l��)�oy��׺���H��E����j#���	���O��q��	}��-�����͵��CU�pk�L�##��]��N�a��.[�}�|�DD�5�������2#�W�X6�!e�&˜|��(�:����%j/6���-�I�S_ �Z͟�<����Q�}�h�~<�XԬb�����d�.7�3�0�0&qk�)�(������Sq�?��i �:^��c�����wi�.�>�E�����o� ,�ɉ\�X�p�pk���yax7�Ԩ����Ȥ�W�|q�������eI�ł�ט
`CzN�k���f����_��|:��S_�?�����B��CO�z��)�r=K�'���6�l;��눅n\^ň2������W;�]��]�{@�QA3~��ہZ���H{_tKT��;�+��U�a7�UQ�"F��kI&�n��6U�Qԡ���L���!����3fvlm��GV���8t�e/���ĭc���K�#�[��l����]%���iB�aBTznH�bQ����H��67�ϯ/QF/�;��fKUN�/@?�5})���AS���n��^���(M1��!c϶o���=t�saGB�]�1�;��&�ɽL�Y �<#���]���\���F|��q����R�B�-���F���� �����v%�nP!��_��61e����ݳ�=fI��y<��^����3]#�a-<�A���M�>�"�D�WJ|�����\q3�~X�$��ݝ)��#M8����"&���7��{i( �Bc��E���ȁ�pP�&"e����ځJuy��2w�U�:�:���vuN���0��|����18L�^~��F⟷��>a��}Z�J��Ehc���+�NM4���U"�,zMir��b��<��KhN�*��z=G�S��Ϩխ�Lg�y��}a�nWѝ�_�ԖG�
���3�(B�X+y���6�!�c�l�e�՗]k!��v��}�㈑C����