XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���8��M؎�h֋1"���ɡ��i@��=ʒ�"ԱP��i� �O�oDp;���'C>��q��|��,���t��.X�������=�p�u�~��Jע�Nk�,d��˜,f��5��C+�j��-�,2^��A�h<��N�&��x���8��p`�}�{��q��O���]���I�Tt��w��r�E-�r��(j`}�{B�����������P%�%���.c[6ņ��S(|�?� /6�7����cF�MU�+�D���:N�gv��|���O,�3��+�JBP��+�U
�Нȶ,����i����+���2?G����J�2Jt��M-Z3�۔��T%��euESC�i!>�G+�ǃ+7<*�	�F�Q�p��1�e��ʼ���2LU����WK:ĎB'����ВP�=��
uM��½G�03>�ӋP�]}H�ls`���嵟#�2�S�gK*I�ԥ��?:�lƂ8SC��Әv�l�t����a�:~���
]槖��c�c����2�N�=�ٶ	ɖ�5f�^�PxN���LK���3���T��S�忢�]Q�ªC�w�:�N��}��}���M)�j��pL���2X�S�,W%�s���<��a)�U��ލ3U6n�4�O���(��.��o��Ys�,@�ٓ`�e��J��hmLi7��(M�����ñ�-~��La�L��ޝq��:�����}O�ur���[[f�O჋�zRp<{�0��O�>�1�T�TL�XlxVHYEB    8625     ee02}�)28]���^72Ŝ6�ck��̕0%�R`0E�W��f*�(0Ơ�\bbQe;b��(ɖe�<<��� 4@��ZS�h{��#8�g7��� `��%��Е|�]/^��<w���+���H�����2�����[��빶��yNj����¡E?����늆�5"r��m��E���Ƒv��?KA��qB��O8;R9�{�]P�6�y�f_�/�E݅�7�FM������g�$W�>�ߗ�%q���S�3]�"��zm��;�i)zB�j�^�ŝ�Z��U�u���} [^��_#1@��sA���x^ϊ��
1+-�=���Q�N��x�Ũ���|<��F�qF���� �Z?��q2�|�)��s�ؽ��m�v4K�vlzM�b�k%i���#���w]Q���pS�87Y��]�#ϙ�Sa�GP�,��������&hXo���al�R�qg��H����;Q&c	�?���J�s��򕲚�[`i�S)��Ǆ�@�Gd3��Ո����8ҁ�9n��!5�������������NW��H�5�8/���=8m��m+���B��#O�D�,{��6�2���"F�\9Vn�3��lP�v����(����vĶ �w�k���\�U<�A�R�~F�ٸ�CvA>J_FSM:M�2.�?v��U�b�^��ݒ'gfr �]�.�?l�,�!W��R�#���� !�p�eT]�x����Bf �Xr[�;�vK5qf������C~?C8�p籜ǁsm�r�r�%��X�эѠq���׬��Lɭ�K����.?�Ώ�t��2N"t�Ԋ4Jp{|��w�Ʋ`Ʃ$��f=1�(��}xb�)q7��w]w�Y��?:��d�Q�W�s�[`�y��I4��7�����4�0*�`��X�(C�9�C!q��*�C�J�0�6U4��g����^VS�qKtj銽P���Y�г���31�[Y������W%�Lp�'	s�C���?*n_6��sIR�p�&�Ik5_���0H.OG�t�&V�d5�X�y�a�u�a|g-��@�m�u��_8m�m=�]et���)_�J�bY:W<'_f �I�δ;T~�<�i��{�W�t�+���M��u���KW����_�}�5y-]�` �'���)��o�����Fҍb�߉��)*{�?Ky���mI(��|{)3���zsU>����<�/Vg7�hF@f����O�U��7.W*i�+�h���맰����Dh@��M=,�`�U=�w\��}`=\���H��OuBg�vݦ���pYep�7���hr>��+ꆜ1vۖ˪��]z���69�<�כ:�|7����u�����2���$�y��%�M���64Z@c�9� �Mk�؆e��&��}�]���};�?mֿ���C�H������U�-t��ވ�<�f��+wEQ���-6�||22)�/e��<�L�;�1��2v��=�;O�<��U�多i�0O��6����tD�N4��Lz�\.B�!��5:R2"6���[.׽"4���H���t�������gF}�ح��Gt�F,5���_�6,�pwrԿ �~U����<�I#F�dqDe��C|F��	�2�H����B�3��n������r���r��B#7�o�$�O�NS�E�LŇ�Ĕw���	��Q7�q�[��O��a!l�[s�����3�T{� t�<��;Ǽ�����<[qcʹ�$�M>8��c 0M<OցQD(��Z�W9���5�:y�*��e	Al�
��CbR��ݔw��t)A�̷�l���0Tg�)�[,�&,")k��y�� �Oճ�)I3G�0�ĝ��9���cDE౑��P�C���J]�z���ڛK1��>�t？�Н�l�ϴ`���!$ ���M������H`�Fvk����c�Z��)8LF�I�o����ΠJ�d���������b�������ǒ~��I>�������;��t�:qO��s��m��\�2А�Te�Q�)c9�}ˆu��u��5�L�5-B��~:������-��v������c�d�v�4v �BEcjC��	%��VC�U0�9%3��1�,�y�����8��K�b���x�d��}��b��/$�AY�uH�M��G�pZ���������kȯ\I��]����s��wp������`�J�����q��D�$m��B���&л�<��4Ix���k���F��Ct�E�����f����px�k�TCR�OWX3a;���+�s����IW*��ΐLaV�'���e=����Pnh���r�μ�/��`.�B�L��ل���K�#�z�2?F-�>J7��4�XN����FP�v��诨�KNH��+��dc�2[P��&7��;��w��&0!�H���$C_����vn�F��$\f��kBY�sF")�
�����Q��G_J�v�sk�Qo��gw���ri��x��Z>�BJ\�nSr�
WG��t��ƚ�,G2��u��w�J�u����9q��<`��zZ��V�$�;�W��Kr˄]Glo���Rtg��O�6ڧmw0]�h�`ͤ�R�J<�`߰Ҳ�"Cw(H/���F�˸��� <:c&*�9�\���cR���Ϯf�x�j^)똈5J��K�!�'.J�ou�FY�TX@���X��|H�q�b� 2�E���Ͱ�M��Qu]c����f���P�}̜��hO�guM��
T���>�X��ڼ�
H�/���8����&�J�?@v��g���=ܾ�m��`���m��ý\��hѦ��ŝ�J�,=�� �p���r���D����#�tDj͸���ͫ��M"XԚ�>M�Tژ8�$ ���i#��a�I�O9
M*���d�Ē����},�_H���%�3��s����� �8mz�W��uR�,@�R���-�a��h�����`�<�C���6��e�z�t�%/1���E1��/߬i��\�VfG@*�*�N�\E�	���10�wU�����S�Uґ��!t�Z4~��.OÇ��"�k�V�c�1X��U��Bထ;_���:��D%z�1P��x��ܛ�G�1���^Mk��������|����h���ʀ�e*LC�1���@E�+6ȫ�o������U׎�wy�oz �TFp��AUy6_�'❀��+�K��<�O�����Α��QPPBb�����_c�E�3����a9�O@�mz T�1�s��Јo��G4���b���@1��>��?z�N�\={��oo�����;�@$���iqd�ŊM��t����Z�*��0��)i��Н�d��@�[�PF��D`g����U����^��DvR�[�������=��}%;{$�$M�N�J�F�ا3zn9R(����̔5���@��œ��;���	�ҧľ�j��]�<��-%?+0x����F
'�F��%�a�,�'�l�5�b��NEQ6��U!O��
���r'��ns��_�!,m���?�8S�闥����YwsHF��8���@�`�G�4ۺ��	�N�|�O��Jt^�~�"�d&�gX��R�67���(�7}�z�~�b�#�P��%Z��A]�M(#P��1*�벫�۝�Eu2m�)��*y��A��+MXR.)�4$I ;^F�'�d�J��p&l��B�9�=	�/��Ui���sRjr�C�4��$N���B]go�q�؍u�`�&�e�(*jj�󌼒�t��d9��E#���K\K���\