XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��՛��*�u�c�c3����v�*��cL���aV�Pp4a����@� {|�`�%]�|Z�4�G�����٘�^t���"9}.�*�|�p����|� ��MĄ
VE���1i	��lY ��?@�*��x�	�1\v���~"�(<�|���W��3�?"���4��Z*������hT���&��+{Y -K�L(7���w�'������2$w�i�=�a&!T\�^
L�Iq����P�C��ҵ�H�6��x�Cz�W%!i�fA~���M?�,?��b���)�5b~=�L��k�C�6gM��4�¿�q�:�T.�5����o�`�ʯ��	�EU2���hM'�9Z�}���`��y�`�&㻆e����:��7��2l��A@����a=��pk��o+K��W���4%;
��S�p��[�S8����L|�����TS�T4� 	������5.��+�~1Ⴍ[���b��A��T��-�N���	AC����(3H�x �|z��&؝�G���'I�b �e�#:<�����<{�:��T_��ae�o�$�D�[�x�
g���Qȃ��6�}�I�����SS	�N��7�{�"����������0b[y�O��q����J�P�������QęxS�a���B�&���a�S~����IKq)*v",�<�X#���<}�	=/��f�N����v�����!|�8�"��vf�4�\^�2�3b�������}qr,�IXlxVHYEB    11e4     520�X�7�2sy"��?'b�fصͳ�L�`��S���C�qSkvYƇ�54n�+v�����^�e��a�Uv���]����9��xK��u�7�t1��c�z��8َ���mD��#�����7L����*����*S�:ff�-�GU-�����Ɉ!WX+N��@���O��qmW�4�H����jpf��jt�ki�r\E���H0��9���i{�P�퉀b1�����.V��"F�LzlƑ�I	_y��,-Z����>L����^��I2���T�����ʼ���q���i�� ~
6S63f��[@D}{X=�gP�Q�}�:*�:-��WEw̾GU�5E�^�y��@�����/���	@�I�\��dH�P�I�x����*&г4��! 8���V}1I�J6Z��%"!�OA!�Bt'픔'u�s������4��#��f���ī�Ph,g��wH��J>�ɨ&��+��³ר�&�d�+���ɵ�o���*�A�SX�*��1~�
�8I����3�uT��Z�4���$3�ȋ�@1�J��G���0h9�( o1��@B�_�}��@�P[{B0����D�uy�W��X)��6�ԥ�oV7Y�%!�n��Dޛ�"�eE<O�8��}jj�Uf�4T"���Q��m���cRt�.t߬Y�9V�Xʦy.�f�v��0T=˶p*�M� a�I72@��5�+ZH��76���]F2X��B%3�W/�ύ�����Ռ�Q,B�H��_a�Jp��W��92Z��#Y�3���>~��<Knfg$������^��^�y��Ml��;�zfc�"��h8��z�vJ�U���=�ß���5֭�� *�H���9~�h���._̡��`��[ �Vk�֢�IC��@��7��e�Uù���9�Xf��1�S��<�mq�e��
"H���UBG�h?����l���H�q�j?�*���n�M�R�:wwM�@���u�l�k{`5�%h�ɒy�;p�ĠNϛ����j��NXY�]�����1�`��6��#�E"��'��hn%��y�u܅��l�;_։�P�Ot��Ϙ��[~�7;�!�����6�.�~cVlIȑW?�ޥ�樳��~}��s<��u���8�@a��2���o�b�[ؼ���DvT�w"�
�xWb�������M��L�ڤ-�?}r��r�$���,n�x ��}[h}��u�GVE��Ѐv����e��'ae$�4->���4?��_�:��py�&�M���FFXӟw�EĔ�n�^��̎��C](����7