XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���=���t�go9-;��݄��=��HF�D<�R3��l]@��g-�������t�ڤѷ��2��x���й�A|]�����P�g@��0֛��1A� ��m�����[?�d��z�cUrb{y1��82$'�hW2�K��"�$6);�
E��yUb�b���R�`J����q^���D���:p�M��"ỷ�
��r|��Z������g�j85�Ex�i(����$l	C.���Vnk�U�9w�6�eM<f1��a�\�E<x�Y�gA�0$m���h]\j���-fu��b.�;eN�E�����X2�f�=D�ÎG/�*g����̬4���?IR��N w����ޚ�u�P'��s�L�����ҡAh�o���T#��l ��Mɹ�@Q�����Hٔ�wwv4�!�"��){��ܕ�]�QDz�l�J�������� ����ޜ�Ej�Ӑ�������-�H�|��X��/���:P[�3"�7�^�e8�Êd�^���������3��_�H��m�S�e��T��.{`R�m�,l�����<�$6N!G(��(����|��ZoP#橅��s�yK��q
y�MS�6~&-��ir)>������,L��$�C(���,�6[	��A�:,kva?�r��<űOq�7։�R��+l��I�&@��7��b]�)����q��E��/e�sꛘ����6������G�V0��H��������,��q^�U/�ש��M]�z�XlxVHYEB     b05     370�	%dj�4k����I��d��e��9���KB�|�Y�!� �6ڱ5�-����XR ��e[{���6:�@}R5�`[��݌Z'����	i&$��B	�<ˈ;�W+h��s5Ɍ�w_�LR�?��b�eO�7�-��N�^����
r4���t��b o��y;R�S�ţ{�-e�Hr½t�ޖ/`{�5��X�=p��\Γ^~��>8Ɂs�=`(�/�:��ƀ����3Qf�c�����4�R(�Ԁ��@wÙ�o��������O��n����9����&�+p���,��3w��[?�T��'jǮ5Z����`�>o��{d?{��	����lv����`n{Qb^�+ߚ�C�LݶJ�&m?�6��/4����+4��}=!�+��Go<���X��E��qWA��R>���δ0@�����c��չ�m�L����!V���J�QJP�E�P��_]���c�$T�r�[=���&'k�D��7�o�C��/�#���v�MF���J]Q:+�:�T��P]#�ɶ~���%r�@:ʏ*Q��޺^�|���TD�#��pqB��ar�*����F����*�f�3������7E`z�1Q�vqK#�y�Q8����Y��k0���Q�x_�d�>$9���N5��j�-�'8��۟_��^�u��µ��]��|�b:�N���*Y�wђ�v��ɤ*?N�S^³I�I��u�Y�2��S:�(��&�� \�vA�� RFT�MOiim>Y�P����e�t:8t�O���������X.j駞|ٱ^P�?_j�!c+ ����C؋�
� �����怗��Џ����ʧ��b�+�
`�}�����2$#�FǍ4��!��j�s�