XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}�+(�٢"w�^_��6*�3?����OB��̚��?
Tl�����dG�:L8؍��фՌ�׋�����c�!�ڝY��p�&�J*���‌;�����%k��yզI�")��{�č�R��p���qRq_'����]�L=ƥ��N������]�m�\`�!h�a�k����A�l�Y�D�K+�:l�f{�0�������R�cꐹ��ӄe���ϧ.�N�e&���ȍ�PG��$V�܀cA�a{�W��&��D������
G���(�s�~He�p�?(� &ñ�U?�-��3Ž��m˫ZJ��	���]�T?4j�e��~!l�6v�G�:�����2�D^/�^oSE��j�,���V���nhS^&��A����%���W���0��M>FX��]FB`��F�de�9\|;s��"s��.5�>�P�L�z>�ɮ�,=gcm9�@X�-�ٖ��ݎ�Ⳏ�+*��R�]��<\�U2�H�
��U~�3|H?�z�a������L����6/fӉ�����@����Y�HVxv�r����>O;Gh��9��85����D}L
��A���Tm�3v�.%	��:5�Ҳ�E��������@��=�W�%w3e|�$*s3�ulWۍ��ه��og$�:��őCe��Ŭ���Q���� �B~�sa����Km���rp݇l}�I��Źg�
�S²����Des���/a��,v���q*��\�J�;5P�.�E��@㺛�e<2e���XlxVHYEB    1d51     7b0H��T2�5���V!�%*n������X�&R�/��V_�s`��J2Qw[h&9��ĕv�?�;��#�N]a�}xS��BD�G��?r�Y �J3K���Dfe���QrOV��J�9n��7�u*���)24��/����s*p�Z�;��rԮi�xH�q/���-��℡���-�Wd��d9�EX,�^�Doe���.��h��VޟN��Yޣ�ʽ(���@�]m���ߑ�_�n��d�����Lqa!�jyjN�,��~�x�G\�eqI:���no�������GyT�rϒ��w/�k��BiY![�h����f[�"w��soР�]B���Eq�o�\Z�ci3��y�$T�(�(���aE��r�Ȅ�F�$ڛ��d� EE0�b�e}��t�6>�_hg,�vn�$�c�4�c���x��Sf�}�O�RTFĊ+�,�!mv�6����yL�\:���B���j]�l�enn�s������*���yp��w�y�o}-6E�$�0`�R# f7NH�i�)��I����:^�e�Z-����D��b��c���ٯq���@k�+򨄔8���m�*4¯�#�/��L^ȹ�)�%�{$����i��BɰJO�c���8�n7�3BgMUHZ�T�ˍ���i�[e:�3H��P)(�B]�oL��3�Nd��èx�߱��DEH��9ͥ�ը��/�v	+��t5� (�\ظ��F��ń�Q����v���^R2T�_�i_��:�B��r��R��Y��V��T��a�%9[2/r&�>1�+؃�4�0�S��sw@�7YZ͌\�����^<~M0�K�?�B_������땡n(Ξ.(���,�C%�`��/�v��6��u�ɗ�4��<��r7����ֳ����~�4�;��~�G�:!�'Km3��_�c�G\���χ��w�J��"]<������%�a)g:��ց|��!�9"S򾦠q��u�4o�`{ THj�p +RP����|�W*�L�i��2���L�&����_h����{NFvP���dQ��*�J�	,!�:}S�g�fΚ$�������6�$�v�X���U#r���Xd�)n�D�
�þ�#\=S����[�l�?\C���?��~>����`��$L�w�|\��LW?��l���$�E�w���#���8;y+��˿�V�#���ȥ�K8�~a�ͷGy�k��]p�@kp����kGo���]��"2L�֊߉�M۱w��R�jܑ�T���[���gY��ƁFãڪ���x�4't�X�b[�d����z���j�"S3ĥ���1ɤu�U@�ɍFS@a�o�[m�+H�Zm��2�G�M���\v�-l(�C���9����t�DT�]St�L�w�lq ��^����S�;���8)�τP�b|��
I��	�� ^]��;KH����K3�Zg�K�]�j��s��hga�zU��'�%;aueM+��J��q��E��:� .������|v>|���$5�j~�B�Q�|�<r=�dh�W�ٚ��h��� ,�R7.��u`=z���NN���c#�(��j�E���w�K�8*�)�K�O����.���\@��8B)4����{�8�Yy{L끵��/]�h�Q�+p{Vj1��A�/}��ҲQX������f/�l�\1l��H�\;Cr��]��m8�|=� wW�}a��AҖ�"��JT]�h��Ӱ6deotPC��Q�<��थ��j[M#�/��m��<���2�ה ԅ���y����!��#����y@���|�(	�C�q���\� ���N�'1X�ޞ��$�3�{VP,��}ۛ#�]x������a`�mI@�B�"p�#�t]����!�3;�~:��)����q�,�G�]r�k��s6?�:��B