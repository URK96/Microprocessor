XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��L缝�^a��,^l�{��
�N!bL��'�g��!��sO����ϯB�Y��@�Ҷ����,�%�P�������wnq�7��G6$���-) �@y�6Z���"��2s9�:Ob�^�v�/�xOy���}vF�tm��ɨ�YB:���"�mt�A=6Q�*���C"μ��0�^]}�3BF��[R?��O|`�0i�Cr�rW6��vD���Bp���U7Z� 1u��1��3��N0-�찼��wӉ0��]ڮ��T�}���̒}�^�i����}�Ok+C�|��]�,>.!c}�K��9�)dP*����ݿ傢9��S�C&gf��9?e�.�bI��ٶ?9I� ݥUO8
��	p �;�u�;�I��IzM\���H��Jy��G}�)<CL���y0h+�֯�3D��\'y_�����sI�*�oAf����?���yg���Vo�T<2}���ܷ�6ArQ�$�
 \c�f�w�0�2�kg����IX���/L�y]
?"���w�,����ur� �˟o��>T����|� A~�5�(E���7�����.i����Vŵ�r�!�bl���?&����$���F	!�łb�In7q[mgy�.��,s�AF�QX�^E��V�E1�.�ÄT\����N)��rPV3���c���y褁Y6�F�L��Q;}�/����/-�e�,�_uq1;�비d���(W_͘G��͗�F�O<�.	���f������a�~^���7��XlxVHYEB    1b22     760�a��z�ܻ��@D�(`�a+}�*^2�C�ų���* �[�F�!�\Va%��c/S�M	�Z^3S٠��O�4�]�<w�gQ�
=܈�D��`J�M��h�P���6�sI)"���T�e!(�c��c��1�5�5^u�Q�Or����U'�w(W;����t�M�ʉ�K�8;����diD|4j������u�w.��k������J;P$jCdCX34!�s�����Yj�Cxv��n�%�8h%b��<LG��y>-C!�
���K���{�[,.�
�p����!��U��y>˝�����x�q�b�q9�X��EJ}n?7��[�J��ܾǻ'��YD������6��u�����z��_��Ϳ_^RA��A�?˂���N�[�	%2�Ńī��1PU��� �,���2�_�w��Э�ݠo���C�{��R������k�D��l�nќ�v�z"S|E��z�h2��a�ʷ��X ��x�Ҵ���D��O�w	.�i������*|�d���\eg���B9a�ݓ����0 �X0��x_���@8K�Ķ�� C3����	���Ù���o����]��}������X��!�� &M��d�P6���:Oq������`��$+6��w�7��aY�>)��~ǝ����"�ր�Bjȷ�N��|��Ĉx�t��2���'�ܾ�I�8�"���emp:�1���P��NX�YA�/�C?X�T2��7�h+'��tW���w�����Ç�㝍��g�Y��GwO_t�8��fgZ��h#�aZ.=ѫT!��:���A�'���a��,e%�����������$ 瞷ڒ �پL��?�)_��ι���%R{��]r2���̘��/����'���R�\�n���I5��'�䓻�ʹDRI���<T���1��^ C����f�޼'٢�p`��.�ק������y����#�j��6s5��ٔ��+�ڋ��q����T6���A��1��e_�Sq�n�uo77�`��J'VL_�V����v\���X��ȕ���!)t
�]F+ ��i����M������|A:�ZӖ�XW`��j�i$x�]醷��F��B��_�* ���X^�79�1a����f��\կ���E�^ed�]j[`���2I�ٲ*���:��Dv�;ew}E
�������d�"fD�"1���?{��<�5�.t��ʆ�������3`��k(\�=��;���������w����y} �1zZcv��=m��������Hx����/U������*��0���Ye����M߄�hFg�9��#���#vG�z^AX
K"fy]8!b��~�P45�z���)%�mT�N�Q�
p�_M��p��^�J��C9�|����{�$�h�����RT74m5Y�M�6�=</XL��g#j5�R{K#(�_^ ��>ދZzK���_��4��lm+����:�m�N��_]*��{�4���F���~va������!:���:1:� o�(��_~�g��˵Npyp4�E#�fL�Q1�C��=���U�ε�z�#�m�N��[z�w��ɂG��.�w�9<�s"&"7c�P���D���_�t�E���T�'���TY��X4�L�{\"s�G/MY��c�e]����î�o#���!c��0Q �Lp���u�� I�"�ͧ��|Yo�n�9h�T7IT�ue=�(#�4���N���<d�7d.r�&��]�ݼP��<e�˓�S�U��pV�=�>����Q��޻b�����+c��̟��taս��b�Zj'b0����/Q�H�Y�Q���:����5�o��>�4�P�9�xV�ɟ
-��L