XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����^�������ln�-��EZ�-�� ��F7�Ņ�GJEo�[X��S�G��+��*<X��u�T��N1���^��<G\[��cm{(��Y�y�t`�L���6h�TN �ڀ,��^]5>OA�U/X�-�I�t��D�p_Pt)\S/���Y&T����ׯ)��O0��;2k ���h�#j�.Ձ�x�g��@O��ga�E3T�Ϊ$���|VR����+�W�,���Wd�TZ������{�zKb��J�?E�@��Aw��u�C�u���[�����G��A��ʦ���rZ���ƥT��sK��Y��. ��[ə�Y�%���y"�6{�Mo<�,yW��D�l�;�v��6d�1��c/��!B����+��bד�#�r|�Aһq�<狔��)�7�VF���y��R�
f���H���xQ��%���z�{���WA��{3�ro	.�d������v�m%��s)ЧċB���F? �����(��fr��C�v�l]��%,En��\���B^��~�-ލqS1P��!f���p����&��&L,��f�u�����^�'��j�q9Z�V&���a���!gw��PZW��с\��J��tϿM����M�N^=�.{�'�)Qr�+C�A��є�^1��Ѝ�P����&���@�w��&n���xH�
w	+<ͭ�8W�W���[e�!L��s|�M���f��Q���H�ח�H��,l���9r@ǭ�`�_�BXlxVHYEB    3c92     910��_�A�Ig >�=v�cG���m��7&e��qp7�ґ��;?�k�ē%i�e�)�0�: E�2q1���l��ʢ�P9��>v�y����3T��k0?@�d+y��D�!�k'�k�
eM��n��1�K�y�7��U ��a�%��#O�~�4��2�'��'m�:�'��H[1��,*���u߇u��I�.U��ZK�8�"ժ�D�!L�Wź���N)����}�k�bv �Pz-̻͘Dd_\4m5k��k�i:�I��*}���XI�%�G��ʢ���P$3�TJڧ�x�M'H��Օ��{����H$���X�2�E,6\	r�Ӑ�ݒuwf�"��Sh�Ԯ�=W�t%�?���=vI����)դ�L���Eu���t1#<3Dn��zʢ-)4��<)���N+���cG���+�6�\K���/�"?]�`��5�Ahk�M0*�ء�oZ����$�1m��q2�dGpa����JB��e��{j Ija.�����9�h�D��j��sjJ��[�],|�?��t�ACڿ�-��ڀ*Om|w���P�ş6 g���sO�\�6��Zs�ΐχ�!N펑G�~�z��ԇ�S��w
?}��g�?�������:>X�%��*џ�G��J�D�R�������ښʊ1@��_d�a��o�@�����ZT�\a���^�=���0�˔+�#0+{���5a��u~@g�z-����E�i�������n��$ �[�,=��rMP��c����B���$�4������O��O�����.t� �m-THب�EE(�$8�i�*I�v���ɫ�V����fo��b��&�)cl"�>fkI&�Бm��LA���Vt.%sgo�'���]���n$�����c��do��H�T�����Wk׆��9E�7��.�V��%8�}�а��0�	��v����!ڙ� J��\_YY,{&Xb!�>Pk��#N����+��!� �B1C����@E'<��@;�z{!� ��,<��j������`�W��H��&U�1��S��Џ�Fcod�=� ��t�"��tP}Ԥ�14*��C�M��rL���$K��J�Q�����r�y�j�=�iiH�ra�q��1Uq8������#��BAGYk������Z>���ޏEj�jB� U�2�bP�f���u�/���XpJ�����0�DaԴ�|���8���D���D��o��B?�
�JG}���՟�ZV��QJ�t�._���~>�t6��>B��a]b/ �^�z���Cg<���$T�k"R*Z��a`�>j*������W����b����R>x[�=�{�ۼkd�l}�.�>b&⤹ӑ4�I�!��fE��S���2��1P2j��.1>�=��v�J8 ��.`�����:��b%R�.����\�Aӽ�QѲ|�lXI�����j����M/Mś֝|�^oEU����G�|{Իʜ7c��/QWf���7VE�4��s �����ˡ:���A��k��[��ڃ�=����co�{O3�
G�f�$
"I��ؾٟ�e��L���]_��ӑ]�g��os�6'�]��?�0�/�ŗ�iQ�
0����H��k��z���xCAM�\)B�>�wA��m��;_������x�o��(93�t����y�����(H��}�#����;��0���d]h��e���A>��X��@g���^`�|���6K_����@�,)v�DAb4c��be�=�����@�S�L��Yƍ��ܓ�vЬ�F�o��0���91���	��+�w��ؗ'�v���7]~V�pr�ĖP�����V$�KS�%���=��Ԓ"�H�Ҩ4,�i*H=�����Bx�,�h��7�z�C#u3��$�֛��ڲ�����\���,���\�g�6�x�"u�5������vr"�;0�w�Ǔž���_�$T'a̾x���k�
�����p�I�d��s��s=�L֦�{�t;�/�9���DX|���fA��>h��^v`U��ӳ�?�#���|;�/y3��Z1"˼%�� ��U5��{ u?F|ty|��&��ŉ>Fnh�tu��'�ü�%h^*�6<�=�zCC�����?�ڪ�NՑ�oqu��<����\�ΰ��g*��.w^y�n���b�l��J�͛�h��cceD��'����yG��W�����	m��%�|��b��HLJe�C�t�-��