XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����$L��U��R�T��K�ȇ�r,7�� ����<�~�z���*�lA�����h��ӈ��K/�~)t%l��X��3J5��b4ؓ*�UOv��8�	��ЮL�;�4p�`am@�'�t"��F��ˇ�-z�1F�bF���"-9�kA�0��7���}���DY�^y�#��,K3\��g�	�jc�Zl���XgV���b�ǂ%����F+��ajް��iX S~�3N�$�
F�1N�w
��V�zV��y ��4�fi�R���b4�R�?!��_C��B�Hn����w�u*��MR;3�����ݷ�ڸU�V:Q4I���� �c��xY�J-@�`|�f��I��|?�����\�ͳ��2jB�Z�Qt���kt��)1.5~R��uXO_�f9�ۑ��F����&��0�kF�A���%��kq�n��K_��~�V
!^L���Hcl5��>���/�HY�3a��&�U�������\�d�͇��w��1*@�������^.� �j1���,���`�*ӰH1)U ��������Rm0w���E�q\?�}�ͫ]N��ǧVf�=C�.Ȓ�tf��5���ǡJ�á88lJ���wP���q�����$*�3�0<�.I/�%�%n���ȸh`v��DZ	Jwh��X_}>�[�kV@�!_���$bg�d�w  b'���+��;o*���mMwʣ_Q�X.��d��U;�_���?C"���L��g����ů���r��DU�XlxVHYEB    3a1b     d40�w�������mh�׋�V*)�S��4�ʏ���@�x[.�YEd �B�l�n�c��n�`��#F��ig����mL�X�{��v6�w�)ݐ@�dGr���1�]Η���j��1��M^0_k�\��_��J��~9h�W9�\��Z������wVW$�*�^nC���$�a��8�{�B*w�r����'��3@��\���*z{8_4��\��G���us֎��0�w|_mQi����aY�Hy&5�]M�M_�Z~eʏ8E4�J�����l������5�r<�HH�/�s����9v��*?�7	V�քE�ܫ��0ŸWK/�Z-��A*��4l�uS�rđۡ6���t' � �<݁���zp�A����M,|�*�&:S��sꢆ
ي4� �!�P�9��um?�s�h�J6�Or|`ӡY����~��`J֏��zw���?~�6O�B��l.8�C�V�I~��6ȥ��J�AR:�:��i��2S3g�ғ�3����a1������(�%K'�-(�}�����;"p��'��즱s?8=����د��Zp��B9�v���'(a���;
e(bo�xW����$����|�a׷令zѳ�
6���E��7>�vAU0��:�>��M;�-�,���`%�.�_�P�8_�U|-uU�V��Q�����QG�n�&��Q�^^Ws{�o�
=ܸ����H�l"�rf�݋{���3{�;߄`o��3C�W���c
_��/:�
����¬ۅx^C/c��W�,�����o�f������^� 7� ci'�J���Ä]3�`}7�Ϧ���p 
>J{j��������>t��_�sv�~,�!s��O�c�'�j5��<F6�����R��{�G�X�y9�//�N���dω��|�h���g�R
YRz���Q������_��Zy�c���Q����zI�zM�H� e��C>"z��U�}��L�ۍ�r�]Y�+D/�8��N)�3T��&,�QjXJ���A�)��=|����J�#�4@���-״iD-��o�d�,P�<�BÎ��sΠ9|Vi�lC��D(��Y}��<+�@��zw4����P��7�'R4:7��49A�!	�g'!�T�y�J�3#��L?�Lۭ�� ����Ĕ�����S�ܷ��#{`k�|R4�|&1<kP��q�)���i������2d�s���_�!8*/�|bԔ.2�wg^RE�m��W�=ƞ�}E۟gj�f��YY��ޑ�8CɄ�Z�y5k$+�_R��
82ژ�y6��5�������yڥ��]�V��罡M���^��Z�����������P4�i!A��tK}f�Q�?�щY�r/ȧěǔ.G���'ަs�U���(.ۯI��(�z;��2G��$I+yw�D����pd "�F_G����B�'�Ԕ��~$��H�V7~���j�.'������ [��j]�l�9ܱ�@!Ҥ���Az
sO�T�#2Q|�~����_z\��Y���5�S�2N���ɉP0\%A�<8@O:]��'"	Z���D�0]�	����-R����D��hw
<`��mʑ��^�`oq�2�p]���1�%���B��4��� R��Ru��m'���S�=vPN�������w�񍵀ݺ��`��z%�$,R
RnG��U����藉�h�`���#���`�:I1<v�>P���[�io�A��X,����t	�'Y>�<t"aPx�|�9�������+$�ʰF�9Y\�:Z�[v�PI�`c�.7��9a����xXg�6?��'D��:��o�cINE����3�@����_~{[_-��"�,�^���U]BS\g%3P'�k�Y���F��{w����˖,����S� 2,;���$h'D�mSh��u�¬�$�(����S(��t�׎��"g.o>H��������޹]�1���x�G�ۥ�0�d3D�y6i�qp���˱����Q:��$q,x���t��~
�����6�ΆI��gw��aw��I4�}N����G�O�f�8^��ۗ�69��a��e'����N�2��]�R�-i�Zc��	��Kh�j ��j�nD �z�듌T�}I8�c�<�(s�|�;w�J�,U{���AFPE\�u���廵R�EG>ChyL��B�}Z��8�2�v�tC9�X��ܬ�.BC̻�a���b�������p.d�m�z��qFe�o7-T|A��
2�75��u�]p�%fy���gm�c���+o9�����iD�To!R��|r��J_Ӵt�F(����a����H���}���dz)��d0��8���ћ�6��eQ�6#�-|WD*2J��p[�$F�t��B��KB&�?z{��@�<�?eƐ���n$#*��]��K�C�0��`�\����B�7�	�yl뇜?��}{A�6�ZI`�x��pٟ����$k�?�8���BG����$���kF��e#�83�g����*5,�c��O���1
mڏ;\"�B�ur'MHp���7jA�tĶc�c��?V�n�5�� �a7��Pd+���	���$^`� �c�l������AK�� o�Sƭ���)�^�IEQ���5�/�����Vl��9'*� �7ޅ��}8}�zW�
2�PJ[T뢟E���3GcӁ�.�y�����/��ݾ����ll��@C��Y~�둁��'�;q�rn�����|�d��G��,���,fαe�~[1�Ȓ[���#0V�>O���&�6'Njf��*�S�Ų{�N`P���UQX8�L_'�uw0���|Z�&� �֨.M@����;��̂'Xܢ�R�Pf�	�9>F�TJ�:��wM�w���be-���໒��U�t�2L_7y?I��:��%!�>�&o��M�ƺBm�cB��p����lt�E=��������C�'+�<B���ט���%k�vwmzNh���Cd�`=-wE��e��;���O�������zG��E�Q���c3��GszQ� �e�ojB1���K��uT2�;j�3s)g�iz�wa�ne���u#U�2��L�LV��s� /v�ȁ䥋�d1��%�ӭ��������]�9�g�*?��Yt�Z�����.	�G'_ev���N���b������N�$[��Ƭ��z�II���3��$u��f�g236		`{�B�M{K�k�D�I��9,�4��E�v<��?)�2�3K_������m�$�eV�N!w�*Q�`S!������{�U��lg;���
M���W)\uz��Zh�S�@T;�