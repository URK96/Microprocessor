XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����#B{�}�FZW=p���i�a~/�0�'ºl�uy�Y@DǢt��3�{Bvm.�p���L�65���:�gI�*(�J�j�$�zc�Ygu���,��~k��&���<P��e%tz��;ޡnb��H�8�cEɸd~�C �mnZ
r{ ��t��HC������=��'��8� �@F� �����sӹ�n�(>���[-Xl����G�~��6g(��/�eU�-�)r�Eh| �n�+��� ii$-}E�9�6��N����b����vd/Vo:��(�=|S�C/c���H��t�')� ���\eb-Pc��!�i��͙oi����^�e;&��S����eVd� ��-�~�����+/R>�����c�����X��.�}��`UM��	����'�W��\7#J��LP����B�"g�{�£*������q�Zo�Wsdh`�^$�����Pm�h]�3R�djs��8�u�.��JD�6�A�Sc�nV�)�Tuν^���ߊd:ZN�D���|&�UO[<��X�l�����I>�1V�'սv���7���5lǙ@��!���m{� td����� �f��)yE�?һ  6Nz�4{�(�����4��k�K�{ӫ�X��4m�TpH��&�w�����鈋R`�6I`c:#��	�e�ץ��b����\t'���f�����w��1\�r>�B��1���h�0�5���J���^XlxVHYEB     9e2     330�4%�)m�5�����$�Œjw�t�)n�N�Ї��ŷĈf��f��Juq����믰���ߋ�rV�s���]�� ^c�bQ��q�c"U�S�`C*�;.��v%��?r�:#2r�J�8|��KwGu7HG_�l[=i(���]!�.��ϱIO�5�o��k���u����jse��D�u`�8��++���Q{�����|3�T��B�ؚ�6-�6K k��ޟ�]�w?sN�Z˿��?.�lp3��m���d�5J=�
�߃����9���q��&�p%�9]ȉ�1³�8����ui���RQͲ�H�8����}���������[�#�Q�Fn��c\���3�����]�Дe�c6}�R�E��n
j�Ie�c��Oc�v���$#h4!ɻXMZ�ds��7�b�oXʠ��/�����c~��8�
֙��}��3cҿ��~�'u�u{i��D���!�rm��et������d!4����2t�+:i"��6v�r��;�P����}!'�12 ����U�!8$���5�L����~�p��W!ފY�(���g�3����̷�D�v��]�<7��Z��#�3�ك�=K�.�V�+�W{�_A_�=e�����b��ʜH���Jn�\�펉I����`�����Q�{��֑���b�*4�#�a��$�q�yxm�P������g<�O/jB�FR���!������$�P�,�>�U�Y��e}'~U�Ha��w�&�'9��^`F�[�Y /#N��Dq��#�.�6Z1�� �Zz��M