XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��7;8����9�������I����˚�1B����eRC�XL�%n�����%gw�q��Я6��Y�ݖ�?Isc�t�vx��:��'alY�@v�fL�?��m:��8B��N\�7i"]��=.oy�P?�7�Տ�y�V��4M�iЭ�&>�U~hb���U��kk�K뺲���5Z��_i��x��z�/��`H�3ȑ�vW��º�OZ��d��Ο�̑i6�e�V���ց?�@p�3IL9rDN���pg@��[��A�8���(���95<�
�'���Sb����F�S��z?>��)2K�����*e����a��6��8�4ʷ���ݪ $�B�JY�����zn�0p�vl��Pi�A���H�x���X���Þ�&Ѩ@��4&�!�x����#��t���AOc��I�����Mcg��>iN�ޔ�ي�g�G]`��Zx�3J�'ܟڽg�?;E$y�
0��/y��Z	4�c�J�09�P��g��L,NG�&i'�+1�]T���\�o#�G oH�V��g������>B�=�%_^Q�&WOҍ�����"r�lN��#�l�޷.�(�Tє����p�����	�w?�9��HNѲ���UU�����F%���-����$�M��5����t�U����.H���jaC5��N;Ñ��7gN˭�kq�.i=�n��<Na��^�&�_�h_}����C�V��.]�^2n�cz���.�fu;8i!h�x�)�GXlxVHYEB    2695     680��v'Do�i�����kP$Z�ل�#/�e@�To�����&꡽����3��`bat���a��~ʵAZZ�U�,.ۿǗKqh��ъ*;^�]U,�`7�6Մ�s�3�zQ�G��y�����~�y)�H��+K��Φ,v_��?�YɐWk	:�0�HY�����:]{����������n���|�6�R5���GV��pN�`D8��G�M�"U��0L�Ǎ��.�l�ĺ�H8�+@^ױ���(�@���z��o�+���+�h�g�����{Ӿ�����ѯt���qw�,l��|(�l#���F�rxl���n��(�k'�ҵ����I9<.7��.����m��޹�N��IR���'�b��°��
�p��~:�!����R��H_C�8��٪� ��y@��`�G����%��K�¥[�Z��Vą��s��)7�I[�솥cR��
|�jRl�ò�@�`g,X��*�d3@�~]*Y!��n`�vdQ
:��f<�wox��]��c4�ǂ�1����(�u�ݬv 
A|���~�@�1�c��p�����"
^����0��f6W��,q�q4.
,��($�;%�@���e��7�ZR�uJs[n
�P:�b�h�W�l�ꊦL�KX�h_�C���*�o�mGg�n���p�&U����D�"��u�¤�O�F}��@QK$�;�[m�m]L�>�A��_���-Q��B��=yI�
�Uo�6����K�_\�����	��Y���]K�f��ܚN�!I��TS�Q+sQZ	rQ[��bj��^�Wcu0����G�]���'Z���)��K���{[%��.���d�]�YXx�m�v���ɗ[?�U�勊/)cm�@AC�}1
_�s�����i��a��d�z�fi
�X
y��M0�\��m7[
?5 �t|�gz���YN���X%�z�T`�:��R��Ӎ�}bbYI�
��,�؎��=��plZ�GpRm@&r��]kw���ml�~��@.E�%��mbJ���hϠJ����R��[�@�]��u3� �˾Sɘ�b�Tə���`��\M����U�x�3sL4�`@A+Q�y��� �r&pD�vz�_%P� ���:��PN�)��0ɖ�M"���L�`�bG�L���z����G��Gf�.��i5�t��S��̰�F��\�Ls
F784�J�v�-�X��૵�ש��߬9�f>����]W�'��91�]��X��x��|
�����ˌ���%S�CA]t�E�����(�q��{�L���~���	i�����V�I�AO	A�f��j�59��Q6B���Z��d���uٹ����U�����$�ч�}��!I_I`$��Y��B�s��t`Crk!�Ώ���**v��&�F�P�z�L�|w\6��Ws����4D�Cz��菹j���ܹڟ�b�B���3�7��k��z\7`�YY�|�%��2����y�Y���LE
���>��?��W����� L(vF�:6#j���6t�pX^�q�<џ��-��;ఞ�m�窓]�&Ky�������ͫ7��~�J��Y���ոK���᚝�h��� X�0��+�#��)3��Q����=��ݴ:��Y�?B��^��{^